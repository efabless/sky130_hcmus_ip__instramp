magic
tech sky130A
magscale 1 2
timestamp 1716789169
<< pwell >>
rect -328 -327 328 327
<< mvnmos >>
rect -100 -69 100 69
<< mvndiff >>
rect -158 57 -100 69
rect -158 -57 -146 57
rect -112 -57 -100 57
rect -158 -69 -100 -57
rect 100 57 158 69
rect 100 -57 112 57
rect 146 -57 158 57
rect 100 -69 158 -57
<< mvndiffc >>
rect -146 -57 -112 57
rect 112 -57 146 57
<< mvpsubdiff >>
rect -292 279 292 291
rect -292 245 -184 279
rect 184 245 292 279
rect -292 233 292 245
rect -292 183 -234 233
rect -292 -183 -280 183
rect -246 -183 -234 183
rect 234 183 292 233
rect -292 -233 -234 -183
rect 234 -183 246 183
rect 280 -183 292 183
rect 234 -233 292 -183
rect -292 -245 292 -233
rect -292 -279 -184 -245
rect 184 -279 292 -245
rect -292 -291 292 -279
<< mvpsubdiffcont >>
rect -184 245 184 279
rect -280 -183 -246 183
rect 246 -183 280 183
rect -184 -279 184 -245
<< poly >>
rect -100 141 100 157
rect -100 107 -84 141
rect 84 107 100 141
rect -100 69 100 107
rect -100 -107 100 -69
rect -100 -141 -84 -107
rect 84 -141 100 -107
rect -100 -157 100 -141
<< polycont >>
rect -84 107 84 141
rect -84 -141 84 -107
<< locali >>
rect -280 245 -184 279
rect 184 245 280 279
rect -280 183 -246 245
rect 246 183 280 245
rect -100 107 -84 141
rect 84 107 100 141
rect -146 57 -112 73
rect -146 -73 -112 -57
rect 112 57 146 73
rect 112 -73 146 -57
rect -100 -141 -84 -107
rect 84 -141 100 -107
rect -280 -245 -246 -183
rect 246 -245 280 -183
rect -280 -279 -184 -245
rect 184 -279 280 -245
<< viali >>
rect -84 107 84 141
rect -146 -57 -112 57
rect 112 -57 146 57
rect -84 -141 84 -107
<< metal1 >>
rect -96 141 96 147
rect -96 107 -84 141
rect 84 107 96 141
rect -96 101 96 107
rect -152 57 -106 69
rect -152 -57 -146 57
rect -112 -57 -106 57
rect -152 -69 -106 -57
rect 106 57 152 69
rect 106 -57 112 57
rect 146 -57 152 57
rect 106 -69 152 -57
rect -96 -107 96 -101
rect -96 -141 -84 -107
rect 84 -141 96 -107
rect -96 -147 96 -141
<< properties >>
string FIXED_BBOX -263 -262 263 262
string gencell sky130_fd_pr__nfet_g5v0d10v5
string library sky130
string parameters w 0.69 l 1.0 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
