* SPICE3 file created from opamp.ext - technology: sky130A

.subckt sky130_fd_pr__res_high_po_0p69_T8KQH6 a_n199_n866# a_n69_n736# a_n69_304#
X0 a_n69_304# a_n69_n736# a_n199_n866# sky130_fd_pr__res_high_po_0p69 l=3.04
C0 a_n69_n736# a_n69_304# 0.0134f
C1 a_n69_n736# a_n199_n866# 0.659f
C2 a_n69_304# a_n199_n866# 0.659f
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_K8DQNF a_n29_n1536# a_229_n1536# a_n229_n1562#
+ w_n487_n1762# a_n287_n1536# a_29_n1562# VSUBS
X0 a_n29_n1536# a_n229_n1562# a_n287_n1536# w_n487_n1762# sky130_fd_pr__pfet_g5v0d10v5 ad=2.17 pd=15.3 as=4.35 ps=30.6 w=15 l=1
X1 a_229_n1536# a_29_n1562# a_n29_n1536# w_n487_n1762# sky130_fd_pr__pfet_g5v0d10v5 ad=4.35 pd=30.6 as=2.17 ps=15.3 w=15 l=1
C0 a_n287_n1536# a_n29_n1536# 0.82f
C1 a_29_n1562# a_n29_n1536# 0.326f
C2 w_n487_n1762# a_n229_n1562# 0.257f
C3 a_229_n1536# a_n29_n1536# 0.82f
C4 a_229_n1536# a_29_n1562# 0.326f
C5 a_n29_n1536# a_n229_n1562# 0.326f
C6 a_n287_n1536# a_n229_n1562# 0.326f
C7 a_n29_n1536# w_n487_n1762# 0.023f
C8 a_29_n1562# a_n229_n1562# 0.0619f
C9 a_n287_n1536# w_n487_n1762# 0.868f
C10 a_29_n1562# w_n487_n1762# 0.257f
C11 a_229_n1536# w_n487_n1762# 0.868f
C12 a_229_n1536# VSUBS 0.733f
C13 a_n29_n1536# VSUBS 0.418f
C14 a_n287_n1536# VSUBS 0.733f
C15 a_29_n1562# VSUBS 0.228f
C16 a_n229_n1562# VSUBS 0.228f
C17 w_n487_n1762# VSUBS 12.4f
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_VYCZE8 a_100_n1681# a_n292_n1841# a_n100_n1707#
+ a_n158_n1681#
X0 a_100_n1681# a_n100_n1707# a_n158_n1681# a_n292_n1841# sky130_fd_pr__nfet_g5v0d10v5 ad=4.78 pd=33.6 as=4.78 ps=33.6 w=16.5 l=1
C0 a_n100_n1707# a_n158_n1681# 0.358f
C1 a_100_n1681# a_n158_n1681# 0.901f
C2 a_100_n1681# a_n100_n1707# 0.358f
C3 a_100_n1681# a_n292_n1841# 1.75f
C4 a_n158_n1681# a_n292_n1841# 1.75f
C5 a_n100_n1707# a_n292_n1841# 0.513f
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_F3SB2X a_n100_n1632# a_100_n1544# a_n292_n1766#
+ a_n158_n1544#
X0 a_100_n1544# a_n100_n1632# a_n158_n1544# a_n292_n1766# sky130_fd_pr__nfet_g5v0d10v5 ad=4.48 pd=31.5 as=4.48 ps=31.5 w=15.4 l=1
C0 a_n100_n1632# a_n158_n1544# 0.335f
C1 a_100_n1544# a_n158_n1544# 0.844f
C2 a_100_n1544# a_n100_n1632# 0.335f
C3 a_100_n1544# a_n292_n1766# 1.64f
C4 a_n158_n1544# a_n292_n1766# 1.64f
C5 a_n100_n1632# a_n292_n1766# 0.743f
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_2HXNYY a_n158_n1900# a_100_n1900# a_n292_n2122#
+ a_n100_n1988#
X0 a_100_n1900# a_n100_n1988# a_n158_n1900# a_n292_n2122# sky130_fd_pr__nfet_g5v0d10v5 ad=5.51 pd=38.6 as=5.51 ps=38.6 w=19 l=1
C0 a_n100_n1988# a_n158_n1900# 0.411f
C1 a_100_n1900# a_n158_n1900# 1.04f
C2 a_100_n1900# a_n100_n1988# 0.411f
C3 a_100_n1900# a_n292_n2122# 2.01f
C4 a_n158_n1900# a_n292_n2122# 2.01f
C5 a_n100_n1988# a_n292_n2122# 0.743f
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_24QKAW a_29_n1997# a_n487_n1997# a_487_n1900#
+ a_n287_n1900# a_n229_n1997# a_n545_n1900# a_n29_n1900# a_287_n1997# w_n745_n2197#
+ a_229_n1900# VSUBS
X0 a_487_n1900# a_287_n1997# a_229_n1900# w_n745_n2197# sky130_fd_pr__pfet_g5v0d10v5 ad=5.51 pd=38.6 as=2.76 ps=19.3 w=19 l=1
X1 a_n287_n1900# a_n487_n1997# a_n545_n1900# w_n745_n2197# sky130_fd_pr__pfet_g5v0d10v5 ad=2.76 pd=19.3 as=5.51 ps=38.6 w=19 l=1
X2 a_n29_n1900# a_n229_n1997# a_n287_n1900# w_n745_n2197# sky130_fd_pr__pfet_g5v0d10v5 ad=2.76 pd=19.3 as=2.76 ps=19.3 w=19 l=1
X3 a_229_n1900# a_29_n1997# a_n29_n1900# w_n745_n2197# sky130_fd_pr__pfet_g5v0d10v5 ad=2.76 pd=19.3 as=2.76 ps=19.3 w=19 l=1
C0 a_29_n1997# a_287_n1997# 0.109f
C1 a_n229_n1997# a_29_n1997# 0.109f
C2 w_n745_n2197# a_n487_n1997# 0.386f
C3 a_n29_n1900# a_29_n1997# 0.411f
C4 a_n29_n1900# a_n229_n1997# 0.411f
C5 a_n287_n1900# a_n229_n1997# 0.411f
C6 a_487_n1900# a_287_n1997# 0.411f
C7 a_229_n1900# a_287_n1997# 0.411f
C8 a_229_n1900# a_29_n1997# 0.411f
C9 a_n287_n1900# a_n29_n1900# 1.04f
C10 a_n545_n1900# a_n287_n1900# 1.04f
C11 a_287_n1997# w_n745_n2197# 0.386f
C12 a_n229_n1997# a_n487_n1997# 0.109f
C13 a_29_n1997# w_n745_n2197# 0.343f
C14 a_n229_n1997# w_n745_n2197# 0.343f
C15 a_229_n1900# a_n29_n1900# 1.04f
C16 a_229_n1900# a_487_n1900# 1.04f
C17 a_n287_n1900# a_n487_n1997# 0.411f
C18 a_n29_n1900# w_n745_n2197# 0.022f
C19 a_n287_n1900# w_n745_n2197# 0.022f
C20 a_n545_n1900# a_n487_n1997# 0.411f
C21 a_n545_n1900# w_n745_n2197# 1.09f
C22 a_487_n1900# w_n745_n2197# 1.09f
C23 a_229_n1900# w_n745_n2197# 0.022f
C24 a_487_n1900# VSUBS 0.925f
C25 a_229_n1900# VSUBS 0.527f
C26 a_n29_n1900# VSUBS 0.527f
C27 a_n287_n1900# VSUBS 0.527f
C28 a_n545_n1900# VSUBS 0.925f
C29 a_287_n1997# VSUBS 0.311f
C30 a_29_n1997# VSUBS 0.288f
C31 a_n229_n1997# VSUBS 0.288f
C32 a_n487_n1997# VSUBS 0.311f
C33 w_n745_n2197# VSUBS 22.5f
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_LB7Y8R a_n100_n157# a_n158_n69# a_n292_n291#
+ a_100_n69#
X0 a_100_n69# a_n100_n157# a_n158_n69# a_n292_n291# sky130_fd_pr__nfet_g5v0d10v5 ad=0.2 pd=1.96 as=0.2 ps=1.96 w=0.69 l=1
C0 a_100_n69# a_n100_n157# 0.0202f
C1 a_n158_n69# a_n100_n157# 0.0202f
C2 a_n158_n69# a_100_n69# 0.0387f
C3 a_100_n69# a_n292_n291# 0.105f
C4 a_n158_n69# a_n292_n291# 0.105f
C5 a_n100_n157# a_n292_n291# 0.683f
.ends

.subckt sky130_fd_pr__cap_mim_m3_1_8DB3RK m3_n876_n730# c1_n836_n690# VSUBS
X0 c1_n836_n690# m3_n876_n730# sky130_fd_pr__cap_mim_m3_1 l=6.9 w=6.9
C0 c1_n836_n690# m3_n876_n730# 4.73f
C1 c1_n836_n690# VSUBS 0.686f
C2 m3_n876_n730# VSUBS 2.42f
.ends

.subckt opamp VDD VSS V1 V2 VOUT
XXR3 VSS m1_4128_540# VOUT sky130_fd_pr__res_high_po_0p69_T8KQH6
XXM1 m1_5053_7611# VDD a_4864_8007# VDD VDD a_4864_8007# VSS sky130_fd_pr__pfet_g5v0d10v5_K8DQNF
XXM2 m1_4306_994# VSS V2 a_4864_8007# sky130_fd_pr__nfet_g5v0d10v5_VYCZE8
XXM3 a_4864_8007# VDD a_4864_8007# VDD VDD a_4864_8007# VSS sky130_fd_pr__pfet_g5v0d10v5_K8DQNF
XXM4 m1_5053_7611# VSS V1 m1_4306_994# sky130_fd_pr__nfet_g5v0d10v5_VYCZE8
XXM5 m1_5284_1188# VSS VSS m1_4306_994# sky130_fd_pr__nfet_g5v0d10v5_F3SB2X
XXM6 VSS VOUT VSS m1_5284_1188# sky130_fd_pr__nfet_g5v0d10v5_2HXNYY
XXM7 m1_5284_1188# m1_5284_1188# VSS VSS sky130_fd_pr__nfet_g5v0d10v5_F3SB2X
XXM8 m1_5053_7611# m1_5053_7611# VDD VOUT m1_5053_7611# VDD VDD m1_5053_7611# VDD
+ VOUT VSS sky130_fd_pr__pfet_g5v0d10v5_24QKAW
XXM9 VDD VDD VSS m1_5284_1188# sky130_fd_pr__nfet_g5v0d10v5_LB7Y8R
XXC1 m1_5053_7611# m1_4128_540# VSS sky130_fd_pr__cap_mim_m3_1_8DB3RK
C0 V2 m1_4128_540# 0.179f
C1 m1_5053_7611# VOUT 7.29f
C2 m1_4306_994# m3_5211_1261# 0.771f
C3 V2 m3_5211_1261# 0.0767f
C4 V1 m1_4128_540# 0.088f
C5 a_4864_8007# m1_4306_994# 0.127f
C6 m1_4128_540# VDD 0.376f
C7 V1 m3_5211_1261# 0.14f
C8 a_4864_8007# V2 0.263f
C9 VDD m3_5211_1261# 0.0192f
C10 V1 a_4864_8007# 0.283f
C11 m1_4128_540# m1_5284_1188# 0.031f
C12 a_4864_8007# VDD 1.96f
C13 m1_5284_1188# m3_5211_1261# 0.446f
C14 m1_4128_540# m1_5053_7611# 0.115f
C15 m1_4128_540# VOUT 0.00888f
C16 a_4864_8007# m1_5284_1188# 0.00623f
C17 m3_5211_1261# m1_5053_7611# 0.0415f
C18 m3_5211_1261# VOUT 0.00865f
C19 a_4864_8007# m1_5053_7611# 1.78f
C20 a_4864_8007# VOUT 0.00842f
C21 V2 m1_4306_994# 0.213f
C22 V1 m1_4306_994# 0.399f
C23 m1_4128_540# m3_5211_1261# 0.0111f
C24 V1 V2 0.16f
C25 m1_4306_994# VDD 0.00701f
C26 V2 VDD 0.00314f
C27 a_4864_8007# m1_4128_540# 0.503f
C28 m1_4306_994# m1_5284_1188# 2.09f
C29 V1 VDD 0.275f
C30 a_4864_8007# m3_5211_1261# 0.0192f
C31 V2 m1_5284_1188# 9.56e-20
C32 m1_4306_994# m1_5053_7611# 0.673f
C33 V1 m1_5284_1188# 0.00363f
C34 V2 m1_5053_7611# 4.01e-19
C35 m1_4306_994# VOUT 0.00433f
C36 VDD m1_5284_1188# 1.67f
C37 V1 m1_5053_7611# 0.143f
C38 V1 VOUT 2.75e-19
C39 VDD m1_5053_7611# 10.4f
C40 VDD VOUT -1.29f
C41 m1_5284_1188# m1_5053_7611# 0.0361f
C42 m1_5284_1188# VOUT 2.28f
C43 m1_4306_994# m1_4128_540# 0.354f
C44 m3_5211_1261# VSS 1.23f **FLOATING
C45 VDD VSS 46.6f
C46 m1_5053_7611# VSS 4.65f
C47 m1_5284_1188# VSS 8.17f
C48 V1 VSS 0.865f
C49 m1_4306_994# VSS 5.55f
C50 V2 VSS 0.848f
C51 a_4864_8007# VSS 4.88f
C52 m1_4128_540# VSS 2.47f
C53 VOUT VSS 4.32f
.ends

