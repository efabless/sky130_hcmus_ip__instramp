magic
tech sky130A
magscale 1 2
timestamp 1718246682
<< nwell >>
rect 3816 9037 5527 9177
rect 3816 8195 5726 9037
rect 3816 4781 3828 8195
<< pwell >>
rect 3879 4489 5061 4682
rect 5062 4489 6956 4682
rect 6221 1221 6322 4489
rect 5002 715 6450 1221
rect 3876 247 6956 436
<< mvnsubdiff >>
rect 3887 9078 5515 9111
rect 3887 8349 3930 9078
rect 5478 8349 5515 9078
rect 3887 8314 5515 8349
<< mvnsubdiffcont >>
rect 3930 8349 5478 9078
<< poly >>
rect 4080 8063 4538 8093
rect 4080 8006 4280 8063
rect 4338 8006 4538 8063
rect 4864 8064 5322 8094
rect 4864 8007 5064 8064
rect 5122 8007 5322 8064
rect 4080 4963 4280 5017
rect 4338 4963 4538 5017
rect 4080 4930 4538 4963
rect 4864 4963 5064 5017
rect 5122 4963 5322 5017
rect 4864 4930 5322 4963
<< locali >>
rect 3900 9078 5609 9098
rect 3900 8349 3930 9078
rect 5478 8935 5609 9078
rect 5478 8349 5605 8935
rect 3900 8283 5605 8349
rect 5615 8883 5622 8937
rect 6888 8883 6895 8930
rect 5615 8880 5756 8883
rect 5615 8797 5747 8880
rect 5615 8283 5756 8797
rect 3900 8270 5756 8283
rect 3900 8145 5612 8270
rect 3900 8139 3920 8145
rect 5483 8106 5612 8145
rect 5615 8106 5756 8270
rect 3919 5007 4068 8011
rect 3917 5003 4068 5007
rect 3917 4880 3925 5003
rect 4061 4880 4068 4893
rect 4550 4880 4853 8011
rect 5334 8010 5474 8011
rect 5483 8010 5756 8106
rect 5334 8004 5756 8010
rect 5334 7998 5603 8004
rect 5358 5075 5603 7998
rect 5615 5075 5756 8004
rect 6237 5112 6272 8797
rect 6754 5076 6895 8883
rect 6783 5075 6895 5076
rect 5358 5011 5612 5075
rect 5334 5010 5612 5011
rect 5334 5002 5505 5010
rect 5334 4884 5473 5002
rect 5486 4914 5505 5002
rect 5602 4914 5612 5010
rect 5486 4860 5612 4914
rect 5615 4893 5622 5075
rect 6888 4894 6895 5075
rect 5615 4890 5745 4893
rect 6754 4883 6895 4894
rect 3905 4567 6350 4578
rect 3905 4530 6366 4567
rect 3905 4438 5124 4530
rect 3905 880 3961 4438
rect 4978 1082 5124 4438
rect 6150 4372 6366 4530
rect 5502 1265 5804 4361
rect 6150 1082 6516 4372
rect 4978 912 6516 1082
rect 4978 882 6166 912
rect 4978 880 5745 882
rect 3905 774 5724 880
rect 3905 406 3961 774
rect 5630 406 5714 774
rect 3905 392 5714 406
rect 6254 564 6516 912
rect 6254 392 6366 564
rect 3905 297 6908 392
<< viali >>
rect 5505 4914 5602 5010
<< metal1 >>
rect 5760 8934 6748 8986
rect 5760 8925 6441 8934
rect 6460 8925 6748 8934
rect 5698 8521 5708 8757
rect 5769 8521 5779 8757
rect 4078 8097 4540 8103
rect 4078 8045 4084 8097
rect 4276 8045 4342 8097
rect 4534 8045 4540 8097
rect 4858 8045 4868 8097
rect 5060 8045 5070 8097
rect 5115 8045 5125 8097
rect 5317 8045 5327 8097
rect 4078 8039 4540 8045
rect 4273 8007 4345 8039
rect 4273 5007 4283 8007
rect 4335 5007 4345 8007
rect 5053 7611 5063 7790
rect 5125 7611 5135 7790
rect 5807 7789 5927 8925
rect 5957 8143 5967 8381
rect 6027 8143 6037 8381
rect 5807 7610 5836 7789
rect 5898 7610 5927 7789
rect 5807 5037 5927 7610
rect 5959 5083 5969 5265
rect 6028 5083 6038 5265
rect 6068 5037 6188 8925
rect 6221 8516 6231 8752
rect 6292 8516 6302 8752
rect 6331 5037 6441 8925
rect 6482 8143 6492 8382
rect 6544 8143 6554 8382
rect 6474 5094 6484 5276
rect 6543 5094 6553 5276
rect 6585 5037 6705 8925
rect 6745 8514 6755 8750
rect 6816 8514 6826 8750
rect 3810 4738 4791 4858
rect 3818 4504 4267 4624
rect 4147 4360 4267 4504
rect 4671 4357 4791 4738
rect 5070 4619 5116 5031
rect 5757 5021 6441 5037
rect 6460 5021 6745 5037
rect 4867 4573 5116 4619
rect 5491 5010 5616 5021
rect 5491 4914 5505 5010
rect 5602 4914 5616 5010
rect 5757 4976 6745 5021
rect 5491 4654 5616 4914
rect 6433 4677 6443 4797
rect 6524 4677 6925 4797
rect 4306 4307 4371 4311
rect 4032 4118 4042 4190
rect 4114 4118 4124 4190
rect 4306 1007 4313 4307
rect 4365 1007 4371 4307
rect 4306 994 4371 1007
rect 4569 1006 4579 4307
rect 4631 1006 4641 4307
rect 4867 4197 4913 4573
rect 5491 4529 6346 4654
rect 5284 4386 5294 4438
rect 5486 4386 5496 4438
rect 5810 4386 5820 4438
rect 6013 4386 6023 4438
rect 5225 4348 5297 4357
rect 5225 1281 5235 4348
rect 5287 1281 5297 4348
rect 5225 1269 5297 1281
rect 5335 1240 5452 4386
rect 5861 1240 5978 4386
rect 6010 1269 6020 4357
rect 6072 1269 6082 4357
rect 5284 1188 5294 1240
rect 5486 1188 5496 1240
rect 5810 1188 5820 1240
rect 6012 1188 6022 1240
rect 6221 1048 6346 4529
rect 5922 923 6346 1048
rect 6572 3799 6692 4442
rect 6725 4035 6735 4274
rect 6800 4035 6810 4274
rect 6572 3693 6589 3799
rect 6675 3693 6692 3799
rect 5922 784 6047 923
rect 5918 738 6047 784
rect 5922 706 6047 738
rect 4128 632 4227 642
rect 4128 550 4138 632
rect 4217 550 4227 632
rect 5419 565 5429 617
rect 5481 565 5491 617
rect 5838 568 6047 706
rect 6083 568 6093 706
rect 6145 568 6155 706
rect 4128 540 4227 550
rect 5922 536 6047 568
rect 5918 511 6047 536
rect 6572 511 6692 3693
rect 6721 568 6731 620
rect 6783 568 6793 620
rect 5918 490 5939 511
<< via1 >>
rect 5708 8521 5769 8757
rect 4084 8045 4276 8097
rect 4342 8045 4534 8097
rect 4868 8045 5060 8097
rect 5125 8045 5317 8097
rect 4283 5007 4335 8007
rect 5063 7611 5125 7790
rect 5967 8143 6027 8381
rect 5836 7610 5898 7789
rect 5969 5083 6028 5265
rect 6231 8516 6292 8752
rect 6492 8143 6544 8382
rect 6484 5094 6543 5276
rect 6755 8514 6816 8750
rect 6443 4677 6524 4797
rect 4042 4118 4114 4190
rect 4313 1007 4365 4307
rect 4579 1006 4631 4307
rect 5294 4386 5486 4438
rect 5820 4386 6013 4438
rect 5235 1281 5287 4348
rect 6020 1269 6072 4357
rect 5294 1188 5486 1240
rect 5820 1188 6012 1240
rect 6735 4035 6800 4274
rect 6589 3693 6675 3799
rect 4138 550 4217 632
rect 5429 565 5481 617
rect 6093 568 6145 706
rect 6731 568 6783 620
<< metal2 >>
rect 5708 8765 5769 8767
rect 5701 8757 6833 8765
rect 5701 8521 5708 8757
rect 5769 8752 6833 8757
rect 5769 8521 6231 8752
rect 5701 8518 6231 8521
rect 5708 8511 5769 8518
rect 6292 8750 6833 8752
rect 6292 8518 6755 8750
rect 6231 8506 6292 8516
rect 6816 8518 6833 8750
rect 6755 8504 6816 8514
rect 6492 8391 6544 8392
rect 5967 8382 6548 8391
rect 5967 8381 6492 8382
rect 6027 8143 6492 8381
rect 6544 8143 6548 8382
rect 5967 8131 6548 8143
rect 4084 8097 5318 8107
rect 4276 8045 4342 8097
rect 4534 8045 4868 8097
rect 5060 8045 5125 8097
rect 5317 8045 5318 8097
rect 4084 8035 5318 8045
rect 4273 8007 4345 8035
rect 4273 5007 4283 8007
rect 4335 5007 4345 8007
rect 5054 7791 5908 7803
rect 5054 7790 5397 7791
rect 5054 7611 5063 7790
rect 5125 7611 5397 7790
rect 5054 7606 5397 7611
rect 5453 7789 5908 7791
rect 5453 7610 5836 7789
rect 5898 7610 5908 7789
rect 5453 7606 5908 7610
rect 5054 7598 5908 7606
rect 5968 5276 6544 5286
rect 5968 5265 6484 5276
rect 5968 5083 5969 5265
rect 6028 5094 6484 5265
rect 6543 5094 6544 5276
rect 6028 5083 6544 5094
rect 5968 5073 6544 5083
rect 4273 4718 4345 5007
rect 4042 4646 4345 4718
rect 6290 4797 6542 5073
rect 6290 4677 6443 4797
rect 6524 4677 6542 4797
rect 4042 4190 4114 4646
rect 5294 4438 6082 4448
rect 5486 4386 5820 4438
rect 6013 4386 6082 4438
rect 5294 4376 6082 4386
rect 6010 4357 6082 4376
rect 4042 4108 4114 4118
rect 4303 4307 4641 4325
rect 4303 1007 4313 4307
rect 4365 1007 4579 4307
rect 4303 1006 4579 1007
rect 4631 2596 4641 4307
rect 5225 2596 5235 4348
rect 4631 2249 5235 2596
rect 4631 1006 4641 2249
rect 5225 1281 5235 2249
rect 5287 1281 5297 4348
rect 5225 1278 5297 1281
rect 6010 1269 6020 4357
rect 6072 3819 6082 4357
rect 6290 4286 6542 4677
rect 6290 4274 6815 4286
rect 6290 4035 6735 4274
rect 6800 4035 6815 4274
rect 6290 4029 6815 4035
rect 6733 4023 6812 4029
rect 6072 3799 6681 3819
rect 6072 3693 6589 3799
rect 6675 3693 6681 3799
rect 6072 3681 6681 3693
rect 6072 1269 6082 3681
rect 6010 1250 6082 1269
rect 5294 1240 6155 1250
rect 5486 1188 5820 1240
rect 6012 1188 6155 1240
rect 5294 1178 6155 1188
rect 4303 991 4641 1006
rect 6083 706 6155 1178
rect 4128 632 4227 642
rect 4128 550 4138 632
rect 4217 550 4227 632
rect 4128 540 4227 550
rect 5429 617 5481 627
rect 5429 527 5481 565
rect 6083 568 6093 706
rect 6145 568 6155 706
rect 6083 557 6155 568
rect 6731 620 6783 630
rect 6731 527 6783 568
rect 5429 475 6783 527
<< via2 >>
rect 5397 7606 5453 7791
rect 4138 550 4217 632
<< metal3 >>
rect 5267 7791 5498 8962
rect 5267 7606 5397 7791
rect 5453 7606 5498 7791
rect 5267 7502 5498 7606
rect 5211 1261 5310 4355
rect 4128 632 4227 642
rect 4128 550 4138 632
rect 4217 550 4227 632
rect 4128 540 4227 550
<< via3 >>
rect 4138 550 4217 632
<< metal4 >>
rect 3926 7582 5226 8882
rect 4138 633 4217 7582
rect 4137 632 4218 633
rect 4137 550 4138 632
rect 4217 550 4218 632
rect 4137 549 4218 550
use sky130_fd_pr__cap_mim_m3_1_8DB3RK  XC1 paramcells
timestamp 1718246682
transform 1 0 4722 0 1 8232
box -876 -730 876 730
use sky130_fd_pr__pfet_g5v0d10v5_K8DQNF  XM1 paramcells
timestamp 1718246682
transform 1 0 5093 0 1 6543
box -487 -1762 487 1762
use sky130_fd_pr__nfet_g5v0d10v5_QXCZXL  XM2 paramcells
timestamp 1718246682
transform 1 0 4207 0 1 2688
box -328 -1877 328 1877
use sky130_fd_pr__pfet_g5v0d10v5_K8DQNF  XM3
timestamp 1718246682
transform 1 0 4309 0 1 6543
box -487 -1762 487 1762
use sky130_fd_pr__nfet_g5v0d10v5_VYCZE8  XM4 paramcells
timestamp 1718246682
transform 1 0 4743 0 1 2688
box -328 -1877 328 1877
use sky130_fd_pr__nfet_g5v0d10v5_9PRBTZ  XM5 paramcells
timestamp 1718246682
transform 1 0 5391 0 1 2814
box -328 -1802 328 1802
use sky130_fd_pr__nfet_g5v0d10v5_2HXNYY  XM6 paramcells
timestamp 1718246682
transform 1 0 6628 0 1 2468
box -328 -2158 328 2158
use sky130_fd_pr__nfet_g5v0d10v5_F3SB2X  XM7 paramcells
timestamp 1718246682
transform 1 0 5926 0 1 2813
box -328 -1802 328 1802
use sky130_fd_pr__pfet_g5v0d10v5_24QKAW  XM8 paramcells
timestamp 1718246682
transform 1 0 6255 0 1 6979
box -745 -2197 745 2197
use sky130_fd_pr__nfet_g5v0d10v5_LB7Y8R  XM9 paramcells
timestamp 1718246682
transform 1 0 5990 0 1 637
box -328 -327 328 327
use sky130_fd_pr__res_high_po_0p69_T8KQH6  XR3 paramcells
timestamp 1718246682
transform 0 1 4778 -1 0 593
box -235 -902 235 902
<< labels >>
rlabel locali 3913 8964 4033 9084 0 VDD
port 1 nsew
flabel metal1 3810 4738 3930 4858 0 FreeSans 800 0 0 0 V1
port 6 nsew
flabel metal1 3818 4504 3938 4624 0 FreeSans 800 0 0 0 V2
port 7 nsew
flabel metal1 6805 4677 6925 4797 0 FreeSans 800 0 0 0 VOUT
port 8 nsew
flabel locali 3912 304 3992 380 0 FreeSans 800 0 0 0 VSS
port 2 nsew
<< end >>
