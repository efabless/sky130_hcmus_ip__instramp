magic
tech sky130A
magscale 1 2
timestamp 1720310800
<< error_s >>
rect -16 -5675 -10 -5669
rect -10 -5681 -4 -5675
rect -10 -5755 -4 -5749
rect -16 -5761 -10 -5755
<< dnwell >>
rect -520 -10586 20480 20584
<< nwell >>
rect -630 20378 20590 20694
rect -630 -10380 -314 20378
rect 20274 -10380 20590 20378
rect -630 -10696 20590 -10380
<< pwell >>
rect 15152 20069 20089 20096
rect 18352 8984 19495 16069
rect 3248 4 19065 4444
rect 16481 -53 20102 -37
rect 49 -1608 20106 -53
rect 9975 -10266 10165 -1608
<< mvpsubdiff >>
rect -879 20025 -771 20049
rect -879 -10571 -771 -10547
<< mvnsubdiff >>
rect -563 20607 20523 20627
rect -563 20573 -483 20607
rect 20443 20573 20523 20607
rect -563 20553 20523 20573
rect -563 20547 -489 20553
rect -563 -10549 -543 20547
rect -509 -10549 -489 20547
rect -563 -10555 -489 -10549
rect 20449 20547 20523 20553
rect 20449 -10549 20469 20547
rect 20503 -10549 20523 20547
rect 20449 -10555 20523 -10549
rect -563 -10575 20523 -10555
rect -563 -10609 -483 -10575
rect 20443 -10609 20523 -10575
rect -563 -10629 20523 -10609
<< mvpsubdiffcont >>
rect -879 -10547 -771 20025
<< mvnsubdiffcont >>
rect -483 20573 20443 20607
rect -543 -10549 -509 20547
rect 20469 -10549 20503 20547
rect -483 -10609 20443 -10575
<< locali >>
rect -567 20607 20523 20627
rect -567 20573 -483 20607
rect 20443 20573 20523 20607
rect -567 20570 20523 20573
rect -567 20547 -84 20570
rect -879 20025 -771 20041
rect -1070 17413 -879 20019
rect -1070 17175 -1049 17413
rect -2378 16332 -2244 16347
rect -2378 16217 -2364 16332
rect -2258 16325 -2244 16332
rect -1711 16325 -1646 16838
rect -2258 16260 -1646 16325
rect -2258 16217 -2244 16260
rect -2378 16166 -2244 16217
rect -1693 14627 -1473 14632
rect -1673 14618 -1625 14627
rect -1591 14618 -1545 14627
rect -1511 14625 -1473 14627
rect -1339 14627 -1224 14632
rect -1339 14625 -1301 14627
rect -1511 14618 -1301 14625
rect -1267 14618 -1224 14627
rect -1691 14593 -1224 14618
rect -1693 14585 -1224 14593
rect -1693 14577 -1664 14585
rect -1691 14538 -1664 14577
rect -1265 14577 -1224 14585
rect -1265 14538 -1238 14577
rect -1691 14520 -1238 14538
rect -2378 13836 -2244 13851
rect -2378 13721 -2364 13836
rect -2258 13829 -2244 13836
rect -1711 13829 -1646 14342
rect -2258 13764 -1646 13829
rect -2258 13721 -2244 13764
rect -2378 13670 -2244 13721
rect -1693 12131 -1473 12136
rect -1673 12122 -1625 12131
rect -1591 12122 -1545 12131
rect -1511 12129 -1473 12131
rect -1339 12131 -1224 12136
rect -1339 12129 -1301 12131
rect -1511 12122 -1301 12129
rect -1267 12122 -1224 12131
rect -1691 12097 -1224 12122
rect -1693 12089 -1224 12097
rect -1693 12081 -1664 12089
rect -1691 12042 -1664 12081
rect -1265 12081 -1224 12089
rect -1265 12042 -1238 12081
rect -1691 12024 -1238 12042
rect -2378 11340 -2244 11355
rect -2378 11225 -2364 11340
rect -2258 11333 -2244 11340
rect -1711 11333 -1646 11846
rect -2258 11268 -1646 11333
rect -2258 11225 -2244 11268
rect -2378 11174 -2244 11225
rect -1693 9635 -1473 9640
rect -1673 9626 -1625 9635
rect -1591 9626 -1545 9635
rect -1511 9633 -1473 9635
rect -1339 9635 -1224 9640
rect -1339 9633 -1301 9635
rect -1511 9626 -1301 9633
rect -1267 9626 -1224 9635
rect -1691 9601 -1224 9626
rect -1693 9593 -1224 9601
rect -1693 9585 -1664 9593
rect -1691 9546 -1664 9585
rect -1265 9585 -1224 9593
rect -1265 9546 -1238 9585
rect -1691 9528 -1238 9546
rect -2378 8844 -2244 8859
rect -2378 8729 -2364 8844
rect -2258 8837 -2244 8844
rect -1711 8837 -1646 9350
rect -2258 8772 -1646 8837
rect -2258 8729 -2244 8772
rect -2378 8678 -2244 8729
rect -1693 7139 -1473 7144
rect -1673 7130 -1625 7139
rect -1591 7130 -1545 7139
rect -1511 7137 -1473 7139
rect -1339 7139 -1224 7144
rect -1339 7137 -1301 7139
rect -1511 7130 -1301 7137
rect -1267 7130 -1224 7139
rect -1691 7105 -1224 7130
rect -1693 7097 -1224 7105
rect -1693 7089 -1664 7097
rect -1691 7050 -1664 7089
rect -1265 7089 -1224 7097
rect -1265 7050 -1238 7089
rect -1691 7032 -1238 7050
rect -2378 6348 -2244 6363
rect -2378 6233 -2364 6348
rect -2258 6341 -2244 6348
rect -1711 6341 -1646 6854
rect -2258 6276 -1646 6341
rect -2258 6233 -2244 6276
rect -2378 6182 -2244 6233
rect -1693 4643 -1473 4648
rect -1673 4634 -1625 4643
rect -1591 4634 -1545 4643
rect -1511 4641 -1473 4643
rect -1339 4643 -1224 4648
rect -1339 4641 -1301 4643
rect -1511 4634 -1301 4641
rect -1267 4634 -1224 4643
rect -1691 4609 -1224 4634
rect -1693 4601 -1224 4609
rect -1693 4593 -1664 4601
rect -1691 4554 -1664 4593
rect -1265 4593 -1224 4601
rect -1265 4554 -1238 4593
rect -1691 4536 -1238 4554
rect -2378 3852 -2244 3867
rect -2378 3737 -2364 3852
rect -2258 3845 -2244 3852
rect -1711 3845 -1646 4358
rect -2258 3780 -1646 3845
rect -2258 3737 -2244 3780
rect -2378 3686 -2244 3737
rect -1693 2147 -1473 2152
rect -1673 2138 -1625 2147
rect -1591 2138 -1545 2147
rect -1511 2145 -1473 2147
rect -1339 2147 -1224 2152
rect -1339 2145 -1301 2147
rect -1511 2138 -1301 2145
rect -1267 2138 -1224 2147
rect -1691 2113 -1224 2138
rect -1693 2105 -1224 2113
rect -1693 2097 -1664 2105
rect -1691 2058 -1664 2097
rect -1265 2097 -1224 2105
rect -1265 2058 -1238 2097
rect -1691 2040 -1238 2058
rect -2378 1356 -2244 1371
rect -2378 1241 -2364 1356
rect -2258 1349 -2244 1356
rect -1711 1349 -1646 1862
rect -2258 1284 -1646 1349
rect -2258 1241 -2244 1284
rect -2378 1190 -2244 1241
rect -1693 -349 -1473 -344
rect -1673 -358 -1625 -349
rect -1591 -358 -1545 -349
rect -1511 -351 -1473 -349
rect -1339 -349 -1224 -344
rect -1339 -351 -1301 -349
rect -1511 -358 -1301 -351
rect -1267 -358 -1224 -349
rect -1691 -383 -1224 -358
rect -1693 -391 -1224 -383
rect -1693 -399 -1664 -391
rect -1691 -438 -1664 -399
rect -1265 -399 -1224 -391
rect -1265 -438 -1238 -399
rect -1691 -456 -1238 -438
rect -2378 -1140 -2244 -1125
rect -2378 -1255 -2364 -1140
rect -2258 -1147 -2244 -1140
rect -1711 -1147 -1646 -634
rect -2258 -1212 -1646 -1147
rect -2258 -1255 -2244 -1212
rect -2378 -1306 -2244 -1255
rect -1693 -2845 -1473 -2840
rect -1673 -2854 -1625 -2845
rect -1591 -2854 -1545 -2845
rect -1511 -2847 -1473 -2845
rect -1339 -2845 -1224 -2840
rect -1339 -2847 -1301 -2845
rect -1511 -2854 -1301 -2847
rect -1267 -2854 -1224 -2845
rect -1691 -2879 -1224 -2854
rect -1693 -2887 -1224 -2879
rect -1693 -2895 -1664 -2887
rect -1691 -2934 -1664 -2895
rect -1265 -2895 -1224 -2887
rect -1265 -2934 -1238 -2895
rect -1691 -2952 -1238 -2934
rect -2378 -3636 -2244 -3621
rect -2378 -3751 -2364 -3636
rect -2258 -3643 -2244 -3636
rect -1711 -3643 -1646 -3130
rect -2258 -3708 -1646 -3643
rect -2258 -3751 -2244 -3708
rect -2378 -3802 -2244 -3751
rect -1693 -5341 -1473 -5336
rect -1673 -5350 -1625 -5341
rect -1591 -5350 -1545 -5341
rect -1511 -5343 -1473 -5341
rect -1339 -5341 -1224 -5336
rect -1339 -5343 -1301 -5341
rect -1511 -5350 -1301 -5343
rect -1267 -5350 -1224 -5341
rect -1691 -5375 -1224 -5350
rect -1693 -5383 -1224 -5375
rect -1693 -5391 -1664 -5383
rect -1691 -5430 -1664 -5391
rect -1265 -5391 -1224 -5383
rect -1265 -5430 -1238 -5391
rect -1691 -5448 -1238 -5430
rect -2378 -6132 -2244 -6117
rect -2378 -6247 -2364 -6132
rect -2258 -6139 -2244 -6132
rect -1711 -6139 -1646 -5626
rect -2258 -6204 -1646 -6139
rect -2258 -6247 -2244 -6204
rect -2378 -6298 -2244 -6247
rect -1693 -7837 -1473 -7832
rect -1673 -7846 -1625 -7837
rect -1591 -7846 -1545 -7837
rect -1511 -7839 -1473 -7837
rect -1339 -7837 -1224 -7832
rect -1339 -7839 -1301 -7837
rect -1511 -7846 -1301 -7839
rect -1267 -7846 -1224 -7837
rect -1691 -7871 -1224 -7846
rect -1693 -7879 -1224 -7871
rect -1693 -7887 -1664 -7879
rect -1691 -7926 -1664 -7887
rect -1265 -7887 -1224 -7879
rect -1265 -7926 -1238 -7887
rect -1691 -7944 -1238 -7926
rect -2378 -8628 -2244 -8613
rect -2378 -8743 -2364 -8628
rect -2258 -8635 -2244 -8628
rect -1711 -8635 -1646 -8223
rect -2258 -8700 -1646 -8635
rect -2258 -8743 -2244 -8700
rect -2378 -8793 -2244 -8743
rect -1691 -10375 -1238 -10342
rect -1691 -10422 -1664 -10375
rect -1265 -10422 -1238 -10375
rect -1070 -10405 -879 17175
rect -1691 -10440 -1238 -10422
rect -879 -10563 -771 -10547
rect -567 -10549 -543 20547
rect -509 20516 -84 20547
rect 20333 20547 20523 20570
rect 20333 20516 20469 20547
rect -509 20489 20469 20516
rect -509 20334 -434 20489
rect -509 -10427 -506 20334
rect -447 -10427 -434 20334
rect -285 20315 20143 20347
rect -285 20204 -240 20315
rect 20105 20204 20143 20315
rect -285 20073 20143 20204
rect -285 334 -256 20073
rect -190 20069 20143 20073
rect 20397 20343 20469 20489
rect -190 9006 -152 20069
rect 4093 19847 4233 20069
rect 19345 19847 19495 20069
rect 4093 19558 19495 19847
rect 4093 18892 4233 19558
rect 13167 19557 19495 19558
rect 4351 19012 19231 19445
rect 19339 18892 19495 19557
rect 4093 18692 19495 18892
rect 4093 18492 4233 18692
rect 19339 18492 19495 18692
rect 4093 18292 19495 18492
rect 4093 18092 4233 18292
rect 19339 18092 19495 18292
rect 4093 17892 19495 18092
rect 4093 17692 4233 17892
rect 19339 17692 19495 17892
rect 4093 17492 19495 17692
rect 4093 17292 4233 17492
rect 19339 17292 19495 17492
rect 4093 17092 19495 17292
rect 4093 16892 4233 17092
rect 19339 16892 19495 17092
rect 4093 16692 19495 16892
rect 2065 16111 3639 16253
rect 2065 15773 2207 16111
rect 3497 15776 3639 16111
rect 4093 16069 4233 16692
rect 4350 16168 19230 16601
rect 19339 16069 19495 16692
rect 4093 16011 19495 16069
rect 4093 15949 4241 16011
rect 2065 15760 2220 15773
rect 2065 14973 2144 15760
rect 2186 14973 2220 15760
rect 2065 14949 2220 14973
rect 3482 15757 3639 15776
rect 3482 14970 3511 15757
rect 3553 14970 3639 15757
rect 3482 14952 3639 14970
rect -53 13228 1057 13392
rect -53 12635 111 13228
rect 893 12635 1057 13228
rect 2065 12645 2207 14949
rect 3497 12654 3639 14952
rect 4094 15400 4241 15949
rect 4354 15496 19234 15928
rect 19345 15400 19495 16011
rect 4094 15200 19495 15400
rect 4094 15000 4241 15200
rect 19345 15000 19495 15200
rect 4094 14800 19495 15000
rect 4094 14600 4241 14800
rect 19345 14600 19495 14800
rect 4094 14400 19495 14600
rect 4094 14200 4241 14400
rect 19345 14200 19495 14400
rect 4094 14000 19495 14200
rect 4094 13800 4241 14000
rect 19345 13800 19495 14000
rect 4094 13600 19495 13800
rect 4094 13400 4241 13600
rect 19345 13400 19495 13600
rect 4094 13200 19495 13400
rect -53 12599 1057 12635
rect -53 12574 1061 12599
rect 4094 12592 4241 13200
rect 4353 12652 19233 13084
rect 19345 12592 19495 13200
rect -53 12441 3623 12574
rect -53 12090 111 12441
rect 893 12435 3623 12441
rect -53 11330 -36 12090
rect 95 11330 111 12090
rect -190 334 -151 9006
rect -53 8998 111 11330
rect 3459 12089 3623 12435
rect 3459 11329 3472 12089
rect 3603 11329 3623 12089
rect 3459 9000 3623 11329
rect 4094 12486 19495 12592
rect 4094 11900 4241 12486
rect 4354 11994 19234 12426
rect 19345 11900 19495 12486
rect 4094 11700 19495 11900
rect 4094 11500 4241 11700
rect 19345 11500 19495 11700
rect 4094 11300 19495 11500
rect 4094 11100 4241 11300
rect 19345 11100 19495 11300
rect 4094 10900 19495 11100
rect 4094 10700 4241 10900
rect 19345 10700 19495 10900
rect 4094 10500 19495 10700
rect 4094 10300 4241 10500
rect 19345 10300 19495 10500
rect 4094 10100 19495 10300
rect 4094 9900 4241 10100
rect 19345 9900 19495 10100
rect 4094 9700 19495 9900
rect 4094 9116 4241 9700
rect 4354 9150 19234 9582
rect 19345 9116 19495 9700
rect 4094 9020 19495 9116
rect 3110 8722 3290 8855
rect 3110 4616 3306 8722
rect 3600 8000 4400 8800
rect 6277 5215 6474 8854
rect 6277 5125 6382 5215
rect 6472 5125 6474 5215
rect 6277 4617 6474 5125
rect 9460 4617 9657 8854
rect 12644 4617 12841 8854
rect 15829 4617 16026 8854
rect 93 4306 19016 4389
rect 93 4243 4513 4306
rect -285 -10214 -151 334
rect 3094 4196 4513 4243
rect 3094 149 3285 4196
rect 3287 149 3405 162
rect 6246 149 6517 4306
rect 9430 149 9701 4306
rect 10718 531 10864 4306
rect 12614 149 12885 4306
rect 15798 149 16069 4306
rect 3094 54 19016 149
rect -90 -3815 43 -27
rect 3094 -130 3285 54
rect 16172 -37 16296 -27
rect 19372 -37 19495 9020
rect 16172 -130 20143 -37
rect 195 -187 20143 -130
rect -90 -3915 -73 -3815
rect 27 -3915 43 -3815
rect -90 -8884 43 -3915
rect -90 -8984 -74 -8884
rect 26 -8984 43 -8884
rect -90 -8998 43 -8984
rect 116 -5114 194 -3642
rect 9940 -3752 10292 -187
rect 15916 -188 20143 -187
rect 10007 -3815 10136 -3800
rect 10007 -3915 10022 -3815
rect 10122 -3915 10136 -3815
rect 116 -5115 9956 -5114
rect 116 -5205 9845 -5115
rect 9935 -5205 9956 -5115
rect 116 -5211 9956 -5205
rect 116 -10160 194 -5211
rect 10007 -8883 10136 -3915
rect 10963 -5021 11093 -4830
rect 20029 -5092 20143 -188
rect 10223 -5115 20143 -5092
rect 10223 -5205 10246 -5115
rect 10336 -5205 20143 -5115
rect 10223 -5232 20143 -5205
rect 10236 -5743 10322 -5355
rect 10007 -8983 10022 -8883
rect 10122 -8983 10136 -8883
rect 10007 -8998 10136 -8983
rect 9933 -10160 10238 -9040
rect 20029 -10160 20143 -5232
rect 116 -10214 20143 -10160
rect -285 -10394 20143 -10214
rect -509 -10491 -434 -10427
rect 20397 -10418 20407 20343
rect 20466 -10418 20469 20343
rect 20397 -10491 20469 -10418
rect -509 -10512 20469 -10491
rect -509 -10549 -82 -10512
rect -567 -10566 -82 -10549
rect 20350 -10549 20469 -10512
rect 20503 -10549 20523 20547
rect 20350 -10566 20523 -10549
rect -567 -10575 20523 -10566
rect -567 -10609 -483 -10575
rect 20443 -10609 20523 -10575
rect -567 -10629 20523 -10609
<< viali >>
rect -1049 17175 -879 17413
rect -879 17175 -800 17413
rect -2364 16217 -2258 16332
rect -1664 14538 -1265 14585
rect -2364 13721 -2258 13836
rect -1664 12042 -1265 12089
rect -2364 11225 -2258 11340
rect -1664 9546 -1265 9593
rect -2364 8729 -2258 8844
rect -1664 7050 -1265 7097
rect -2364 6233 -2258 6348
rect -1664 4554 -1265 4601
rect -2364 3737 -2258 3852
rect -1664 2058 -1265 2105
rect -2364 1241 -2258 1356
rect -1664 -438 -1265 -391
rect -2364 -1255 -2258 -1140
rect -1664 -2934 -1265 -2887
rect -2364 -3751 -2258 -3636
rect -1664 -5430 -1265 -5383
rect -2364 -6247 -2258 -6132
rect -1664 -7926 -1265 -7879
rect -2364 -8743 -2258 -8628
rect -1664 -10422 -1265 -10375
rect -84 20516 20333 20570
rect -506 -10427 -447 20334
rect -240 20204 20105 20315
rect -256 334 -190 20073
rect 2144 14973 2186 15760
rect 3511 14970 3553 15757
rect -36 11330 95 12090
rect 3472 11329 3603 12089
rect -73 -3915 27 -3815
rect -74 -8984 26 -8884
rect 10022 -3915 10122 -3815
rect 9845 -5205 9935 -5115
rect 10246 -5205 10336 -5115
rect 10022 -8983 10122 -8883
rect 20407 -10418 20466 20343
rect -82 -10566 20350 -10512
<< metal1 >>
rect -567 20570 20523 20627
rect -567 20516 -84 20570
rect 20333 20516 20523 20570
rect -567 20489 20523 20516
rect -567 20334 -434 20489
rect -2183 17909 -2023 17940
rect -2183 17608 -2023 17631
rect -2707 17433 -2559 17449
rect -2707 17023 -2559 17154
rect -2695 -10404 -2580 17023
rect -2378 16466 -2244 16480
rect -2378 16332 -2244 16410
rect -2378 16217 -2364 16332
rect -2258 16217 -2244 16332
rect -2378 16201 -2244 16217
rect -2378 13970 -2244 13984
rect -2378 13836 -2244 13914
rect -2378 13721 -2364 13836
rect -2258 13721 -2244 13836
rect -2378 13705 -2244 13721
rect -2378 11474 -2244 11488
rect -2378 11340 -2244 11418
rect -2378 11225 -2364 11340
rect -2258 11225 -2244 11340
rect -2378 11209 -2244 11225
rect -2378 8978 -2244 8992
rect -2378 8844 -2244 8922
rect -2378 8729 -2364 8844
rect -2258 8729 -2244 8844
rect -2378 8713 -2244 8729
rect -2378 6482 -2244 6496
rect -2378 6348 -2244 6426
rect -2378 6233 -2364 6348
rect -2258 6233 -2244 6348
rect -2378 6217 -2244 6233
rect -2378 3986 -2244 4000
rect -2378 3852 -2244 3930
rect -2378 3737 -2364 3852
rect -2258 3737 -2244 3852
rect -2378 3721 -2244 3737
rect -2378 1490 -2244 1504
rect -2378 1356 -2244 1434
rect -2378 1241 -2364 1356
rect -2258 1241 -2244 1356
rect -2378 1225 -2244 1241
rect -2378 -1006 -2244 -992
rect -2378 -1140 -2244 -1062
rect -2378 -1255 -2364 -1140
rect -2258 -1255 -2244 -1140
rect -2378 -1271 -2244 -1255
rect -2378 -3502 -2244 -3488
rect -2378 -3636 -2244 -3558
rect -2378 -3751 -2364 -3636
rect -2258 -3751 -2244 -3636
rect -2378 -3767 -2244 -3751
rect -2378 -5998 -2244 -5984
rect -2378 -6132 -2244 -6054
rect -2378 -6247 -2364 -6132
rect -2258 -6247 -2244 -6132
rect -2378 -6263 -2244 -6247
rect -2378 -8494 -2244 -8480
rect -2378 -8628 -2244 -8550
rect -2378 -8743 -2364 -8628
rect -2258 -8743 -2244 -8628
rect -2378 -8759 -2244 -8743
rect -2080 -9426 -2023 17608
rect -1995 17046 -1745 17947
rect -1181 17433 -1033 17451
rect -1033 17413 -770 17433
rect -800 17175 -770 17413
rect -1033 17155 -770 17175
rect -1977 6914 -1771 17046
rect -1181 17034 -1033 17154
rect -1691 14601 -1238 14618
rect -1691 14507 -1675 14601
rect -1260 14507 -1238 14601
rect -1691 14492 -1238 14507
rect -1691 12105 -1238 12122
rect -1691 12011 -1675 12105
rect -1260 12011 -1238 12105
rect -1691 11996 -1238 12011
rect -1691 9609 -1238 9626
rect -1691 9515 -1675 9609
rect -1260 9515 -1238 9609
rect -1691 9500 -1238 9515
rect -1691 7113 -1238 7130
rect -1691 7019 -1675 7113
rect -1260 7019 -1238 7113
rect -1691 7004 -1238 7019
rect -1987 6896 -1744 6914
rect -1987 5851 -1971 6896
rect -1769 5851 -1744 6896
rect -1987 5826 -1744 5851
rect -1977 -10393 -1771 5826
rect -1691 4617 -1238 4634
rect -1691 4523 -1675 4617
rect -1260 4523 -1238 4617
rect -1691 4508 -1238 4523
rect -1691 2121 -1238 2138
rect -1691 2027 -1675 2121
rect -1260 2027 -1238 2121
rect -1691 2012 -1238 2027
rect -1691 -375 -1238 -358
rect -1691 -469 -1675 -375
rect -1260 -469 -1238 -375
rect -1691 -484 -1238 -469
rect -1691 -2871 -1238 -2854
rect -1691 -2965 -1675 -2871
rect -1260 -2965 -1238 -2871
rect -1691 -2980 -1238 -2965
rect -1691 -5367 -1238 -5350
rect -1691 -5461 -1675 -5367
rect -1260 -5461 -1238 -5367
rect -1691 -5476 -1238 -5461
rect -1691 -7863 -1238 -7846
rect -1691 -7957 -1675 -7863
rect -1260 -7957 -1238 -7863
rect -1691 -7972 -1238 -7957
rect -1691 -10359 -1238 -10342
rect -1691 -10453 -1675 -10359
rect -1260 -10453 -1238 -10359
rect -1160 -10399 -1054 17034
rect -1691 -10468 -1238 -10453
rect -567 -10427 -506 20334
rect -447 -8868 -434 20334
rect -313 20315 20138 20344
rect -313 20204 -240 20315
rect 20105 20204 20138 20315
rect -313 20165 20138 20204
rect 20397 20343 20523 20489
rect -313 20073 -94 20165
rect -313 15783 -256 20073
rect -190 15783 -94 20073
rect 4351 19437 19231 19445
rect 4351 19020 19052 19437
rect 19158 19020 19231 19437
rect 4351 19012 19231 19020
rect 4361 16596 19230 16601
rect 2401 16331 3287 16335
rect 2401 16260 2421 16331
rect 2717 16260 3287 16331
rect 2401 16254 3287 16260
rect 2415 15983 2496 16254
rect 3206 15987 3287 16254
rect 4361 16176 16610 16596
rect 16859 16176 19230 16596
rect 4361 16168 19230 16176
rect 2415 15979 2501 15983
rect -134 14936 -94 15783
rect 2117 15763 2220 15773
rect 2117 14970 2131 15763
rect 2210 14970 2220 15763
rect 2117 14949 2220 14970
rect -313 3403 -256 14936
rect -315 3381 -256 3403
rect -190 3403 -94 14936
rect 2288 14827 2381 14855
rect 177 13010 283 13020
rect 177 12835 197 13010
rect 260 12835 283 13010
rect 177 12819 283 12835
rect 328 12781 404 13099
rect 441 13010 547 13023
rect 441 12835 464 13010
rect 527 12835 547 13010
rect 441 12781 547 12835
rect 586 12781 662 13099
rect 698 13010 804 13027
rect 698 12835 718 13010
rect 781 12835 804 13010
rect 2288 12911 2301 14827
rect 2369 12911 2381 14827
rect 2288 12882 2381 12911
rect 698 12826 804 12835
rect 2433 12784 2501 15979
rect 2554 12841 2629 14841
rect 267 12735 717 12781
rect 328 12572 404 12735
rect 586 12572 662 12735
rect 2679 12709 2747 15972
rect 2807 15895 2900 15911
rect 2807 12890 2828 15895
rect 2884 12890 2900 15895
rect 2807 12864 2900 12890
rect 2953 12913 3021 15979
rect 3070 12913 3145 14830
rect 2953 12843 3145 12913
rect 2953 12791 3021 12843
rect 3070 12841 3145 12843
rect 2952 12780 3021 12791
rect 2952 12709 3020 12780
rect 3202 12777 3270 15976
rect 4354 15917 18234 15928
rect 3482 15757 3585 15776
rect 3482 15755 3511 15757
rect 3553 15755 3585 15757
rect 3482 14962 3490 15755
rect 3569 14962 3585 15755
rect 4354 15505 15881 15917
rect 15982 15505 18234 15917
rect 4354 15496 18234 15505
rect 3482 14952 3585 14962
rect 3319 14825 3412 14853
rect 3319 12909 3332 14825
rect 3400 12909 3412 14825
rect 3319 12880 3412 12909
rect 4353 13073 18233 13084
rect 2679 12641 3020 12709
rect 4353 12660 12639 13073
rect 12881 12660 18233 13073
rect 4353 12652 18233 12660
rect 328 12535 3240 12572
rect 328 12473 3242 12535
rect -53 12090 116 12108
rect 210 12092 216 12138
rect 250 12092 256 12138
rect -53 11330 -36 12090
rect 95 11330 116 12090
rect -53 11311 116 11330
rect 191 12084 273 12092
rect 191 10324 197 12084
rect 268 10324 273 12084
rect 191 9347 273 10324
rect 210 9332 216 9347
rect 250 9332 256 9347
rect 328 9154 404 12473
rect 449 11152 531 12092
rect 449 9380 455 11152
rect 526 9380 531 11152
rect 449 9347 531 9380
rect 586 9154 662 12473
rect 726 12092 732 12120
rect 766 12092 772 12120
rect 707 12084 789 12092
rect 707 10324 713 12084
rect 784 10324 789 12084
rect 707 9361 789 10324
rect 844 9154 920 12473
rect 984 12092 990 12120
rect 1024 12092 1030 12120
rect 965 11152 1047 12092
rect 965 9380 971 11152
rect 1042 9380 1047 11152
rect 965 9361 1047 9380
rect 1102 9154 1178 12473
rect 1242 12092 1248 12120
rect 1282 12092 1288 12120
rect 1223 12084 1305 12092
rect 1223 10324 1229 12084
rect 1300 10324 1305 12084
rect 1223 9361 1305 10324
rect 1360 9154 1436 12473
rect 1500 12092 1506 12120
rect 1540 12092 1546 12120
rect 1481 11152 1563 12092
rect 1481 9380 1487 11152
rect 1558 9380 1563 11152
rect 1481 9361 1563 9380
rect 1618 9154 1694 12473
rect 1758 12092 1764 12120
rect 1798 12092 1804 12120
rect 1739 12084 1821 12092
rect 1739 10324 1745 12084
rect 1816 10324 1821 12084
rect 1739 9361 1821 10324
rect 1876 9154 1952 12473
rect 2016 12092 2022 12120
rect 2056 12092 2062 12120
rect 1997 11152 2079 12092
rect 1997 9380 2003 11152
rect 2074 9380 2079 11152
rect 1997 9361 2079 9380
rect 2134 9154 2210 12473
rect 2274 12092 2280 12120
rect 2314 12092 2320 12120
rect 2255 12084 2337 12092
rect 2255 10324 2261 12084
rect 2332 10324 2337 12084
rect 2255 9361 2337 10324
rect 2392 9154 2468 12473
rect 2532 12092 2538 12120
rect 2572 12092 2578 12120
rect 2513 11152 2595 12092
rect 2513 9380 2519 11152
rect 2590 9380 2595 11152
rect 2513 9361 2595 9380
rect 2650 9154 2726 12473
rect 2790 12092 2796 12120
rect 2830 12092 2836 12120
rect 2771 12084 2853 12092
rect 2771 10324 2777 12084
rect 2848 10324 2853 12084
rect 2771 9361 2853 10324
rect 2908 9154 2984 12473
rect 3048 12092 3054 12120
rect 3088 12092 3094 12120
rect 3029 11152 3111 12092
rect 3029 9380 3035 11152
rect 3106 9380 3111 11152
rect 3029 9361 3111 9380
rect 3166 9154 3242 12473
rect 3306 12092 3312 12120
rect 3346 12092 3352 12120
rect 3287 12084 3369 12092
rect 3287 10324 3293 12084
rect 3364 10324 3369 12084
rect 3455 12089 3624 12107
rect 3455 11329 3472 12089
rect 3603 11329 3624 12089
rect 4354 11994 18234 12426
rect 3455 11310 3624 11329
rect 3287 9361 3369 10324
rect 8049 9765 8169 11994
rect 8049 9675 8065 9765
rect 8155 9675 8169 9765
rect 8049 9660 8169 9675
rect 4354 9150 18234 9582
rect 4866 5015 4986 9150
rect 8049 9075 8169 9090
rect 8049 8985 8065 9075
rect 8155 8985 8169 9075
rect 4866 4935 4886 5015
rect 4966 4935 4986 5015
rect 4866 4924 4986 4935
rect 6366 5215 6486 5230
rect 6366 5125 6382 5215
rect 6472 5125 6486 5215
rect -44 4615 76 4621
rect 76 4495 119 4615
rect 3164 4495 3182 4615
rect 6366 4495 6486 5125
rect 8049 5080 8169 8985
rect 8049 5000 8070 5080
rect 8150 5000 8169 5080
rect 8049 4990 8169 5000
rect 15872 9078 15992 9090
rect 15872 8978 15882 9078
rect 15982 8978 15992 9078
rect 15872 4801 15992 8978
rect 20397 6918 20407 20343
rect 19861 6891 20407 6918
rect 19861 5867 19896 6891
rect 20144 5867 20407 6891
rect 19861 5839 20407 5867
rect 15872 4701 15881 4801
rect 15981 4701 15992 4801
rect 15872 4690 15992 4701
rect 16750 5280 16870 5290
rect 16750 5180 16760 5280
rect 16860 5180 16870 5280
rect 16750 4495 16870 5180
rect 19491 5280 19924 5290
rect 19491 5180 19500 5280
rect 19914 5180 19924 5280
rect -44 4489 76 4495
rect -50 4260 -44 4380
rect 76 4260 82 4380
rect -190 3381 4 3403
rect -315 2478 -297 3381
rect -21 2478 4 3381
rect -315 2453 -256 2478
rect -313 334 -256 2453
rect -190 2453 4 2478
rect -190 334 -134 2453
rect -313 284 -134 334
rect 3190 192 3310 4381
rect 6109 446 6264 4125
rect 4730 405 4880 409
rect 4730 395 4764 405
rect -256 72 3310 192
rect 4730 297 4764 302
rect 4787 297 4880 405
rect 6109 377 6333 446
rect 6093 325 6180 377
rect 6317 325 6333 377
rect -256 -4622 -136 72
rect 4730 -339 4880 297
rect 6209 -359 6333 325
rect 6376 -27 6496 4384
rect 15926 4370 16046 4381
rect 15926 4270 15937 4370
rect 16037 4270 16046 4370
rect 9290 548 9445 4125
rect 9290 495 9358 548
rect 9430 495 9445 548
rect 10411 -27 10531 4234
rect 13593 151 13713 4234
rect 13593 20 13604 151
rect 13703 20 13713 151
rect 13593 10 13713 20
rect 6376 -147 6496 -139
rect 9695 -147 10531 -27
rect 15926 -18 16046 4270
rect 17195 374 17616 409
rect 17195 322 17213 374
rect 17493 322 17616 374
rect 18839 377 19051 4125
rect 18839 325 18930 377
rect 19040 325 19051 377
rect 19491 360 19924 5180
rect 19491 334 19925 360
rect 15926 -35 16207 -18
rect 15926 -125 16101 -35
rect 16181 -125 16207 -35
rect 15926 -138 16207 -125
rect 16086 -140 16206 -138
rect 9695 -338 9815 -147
rect 17195 -293 17616 322
rect 19491 214 20214 334
rect 13995 -314 14416 -309
rect 5970 -3603 6123 -3580
rect 3523 -3642 3645 -3617
rect 3523 -3722 3546 -3642
rect 3626 -3722 3645 -3642
rect 121 -4038 140 -3958
rect 121 -4146 140 -4066
rect 121 -4254 140 -4174
rect 121 -4362 140 -4282
rect 121 -4470 140 -4390
rect -256 -4702 -10 -4622
rect 3523 -5132 3645 -3722
rect 5970 -3723 5987 -3603
rect 6107 -3723 6123 -3603
rect 3523 -5212 3547 -5132
rect 3627 -5212 3645 -5132
rect 3523 -5229 3645 -5212
rect 5970 -5563 6123 -3723
rect 16080 -3610 16200 -3600
rect 16080 -3710 16090 -3610
rect 16190 -3710 16200 -3610
rect 16080 -4613 16200 -3710
rect 16080 -4713 16090 -4613
rect 16190 -4713 16200 -4613
rect 16080 -4720 16200 -4713
rect 9830 -5115 9950 -5100
rect 9830 -5205 9845 -5115
rect 9935 -5205 9950 -5115
rect 9830 -5220 9950 -5205
rect 10223 -5115 10363 -5092
rect 10223 -5205 10246 -5115
rect 10336 -5205 10363 -5115
rect 10223 -5232 10363 -5205
rect 10223 -5463 10569 -5334
rect 10223 -5613 10245 -5463
rect -102 -5755 -90 -5675
rect 10223 -5756 10569 -5613
rect 41 -6580 62 -6500
rect 267 -6506 11093 -6500
rect 267 -6573 10970 -6506
rect 11087 -6573 11093 -6506
rect 267 -6580 11093 -6573
rect 41 -6720 62 -6640
rect 267 -6646 11735 -6640
rect 267 -6713 11612 -6646
rect 11729 -6713 11735 -6646
rect 267 -6720 11735 -6713
rect 41 -6860 62 -6780
rect 267 -6787 12627 -6780
rect 267 -6854 12504 -6787
rect 12621 -6854 12627 -6787
rect 267 -6860 12627 -6854
rect 41 -7000 62 -6920
rect 267 -6926 14043 -6920
rect 267 -6993 13920 -6926
rect 14037 -6993 14043 -6926
rect 267 -7000 14043 -6993
rect 41 -7140 62 -7060
rect 267 -7067 16486 -7060
rect 267 -7134 16363 -7067
rect 16480 -7134 16486 -7067
rect 267 -7140 16486 -7134
rect 866 -8705 996 -8690
rect 866 -8805 880 -8705
rect 980 -8805 996 -8705
rect -447 -8884 147 -8868
rect -447 -8984 -74 -8884
rect 26 -8984 147 -8884
rect -447 -8998 147 -8984
rect -447 -10427 -434 -8998
rect -90 -9106 -10 -9026
rect 866 -9106 996 -8805
rect 1508 -8705 1638 -8690
rect 1508 -8805 1521 -8705
rect 1621 -8805 1638 -8705
rect 1508 -9030 1638 -8805
rect 2400 -8705 2530 -8690
rect 2400 -8805 2415 -8705
rect 2515 -8805 2530 -8705
rect 2400 -9060 2530 -8805
rect 3523 -8717 3646 -8707
rect 3523 -8817 3536 -8717
rect 3636 -8817 3646 -8717
rect -90 -9214 -10 -9134
rect -90 -9322 -10 -9242
rect -90 -9430 -10 -9350
rect -90 -9538 -10 -9458
rect 3523 -9697 3646 -8817
rect 3816 -8719 3946 -8707
rect 3816 -8819 3832 -8719
rect 3932 -8819 3946 -8719
rect 3816 -9007 3946 -8819
rect 6259 -8719 6389 -8710
rect 6259 -8819 6275 -8719
rect 6375 -8819 6389 -8719
rect 6259 -9006 6389 -8819
rect 3523 -9767 3550 -9697
rect 3620 -9767 3646 -9697
rect 20094 -9700 20214 214
rect 20094 -9760 20101 -9700
rect 20207 -9760 20214 -9700
rect 20094 -9766 20214 -9760
rect 3523 -9787 3646 -9767
rect -567 -10491 -434 -10427
rect 20397 -10418 20407 5839
rect 20466 -10418 20523 20343
rect 20397 -10491 20523 -10418
rect -567 -10512 20523 -10491
rect -567 -10566 -82 -10512
rect 20350 -10566 20523 -10512
rect -567 -10629 20523 -10566
<< via1 >>
rect -2183 17631 -2023 17909
rect -2707 17154 -2559 17433
rect -2378 16410 -2244 16466
rect -2378 13914 -2244 13970
rect -2378 11418 -2244 11474
rect -2378 8922 -2244 8978
rect -2378 6426 -2244 6482
rect -2378 3930 -2244 3986
rect -2378 1434 -2244 1490
rect -2378 -1062 -2244 -1006
rect -2378 -3558 -2244 -3502
rect -2378 -6054 -2244 -5998
rect -2378 -8550 -2244 -8494
rect -1181 17413 -1033 17433
rect -1181 17175 -1049 17413
rect -1049 17175 -1033 17413
rect -1181 17154 -1033 17175
rect -1675 14585 -1260 14601
rect -1675 14538 -1664 14585
rect -1664 14538 -1265 14585
rect -1265 14538 -1260 14585
rect -1675 14507 -1260 14538
rect -1675 12089 -1260 12105
rect -1675 12042 -1664 12089
rect -1664 12042 -1265 12089
rect -1265 12042 -1260 12089
rect -1675 12011 -1260 12042
rect -1675 9593 -1260 9609
rect -1675 9546 -1664 9593
rect -1664 9546 -1265 9593
rect -1265 9546 -1260 9593
rect -1675 9515 -1260 9546
rect -1675 7097 -1260 7113
rect -1675 7050 -1664 7097
rect -1664 7050 -1265 7097
rect -1265 7050 -1260 7097
rect -1675 7019 -1260 7050
rect -1971 5851 -1769 6896
rect -1675 4601 -1260 4617
rect -1675 4554 -1664 4601
rect -1664 4554 -1265 4601
rect -1265 4554 -1260 4601
rect -1675 4523 -1260 4554
rect -1675 2105 -1260 2121
rect -1675 2058 -1664 2105
rect -1664 2058 -1265 2105
rect -1265 2058 -1260 2105
rect -1675 2027 -1260 2058
rect -1675 -391 -1260 -375
rect -1675 -438 -1664 -391
rect -1664 -438 -1265 -391
rect -1265 -438 -1260 -391
rect -1675 -469 -1260 -438
rect -1675 -2887 -1260 -2871
rect -1675 -2934 -1664 -2887
rect -1664 -2934 -1265 -2887
rect -1265 -2934 -1260 -2887
rect -1675 -2965 -1260 -2934
rect -1675 -5383 -1260 -5367
rect -1675 -5430 -1664 -5383
rect -1664 -5430 -1265 -5383
rect -1265 -5430 -1260 -5383
rect -1675 -5461 -1260 -5430
rect -1675 -7879 -1260 -7863
rect -1675 -7926 -1664 -7879
rect -1664 -7926 -1265 -7879
rect -1265 -7926 -1260 -7879
rect -1675 -7957 -1260 -7926
rect -1675 -10375 -1260 -10359
rect -1675 -10422 -1664 -10375
rect -1664 -10422 -1265 -10375
rect -1265 -10422 -1260 -10375
rect -1675 -10453 -1260 -10422
rect 19052 19020 19158 19437
rect 2421 16260 2717 16331
rect 16610 16176 16859 16596
rect -313 14936 -256 15783
rect -256 14936 -190 15783
rect -190 14936 -134 15783
rect 2131 15760 2210 15763
rect 2131 14973 2144 15760
rect 2144 14973 2186 15760
rect 2186 14973 2210 15760
rect 2131 14970 2210 14973
rect 197 12835 260 13010
rect 464 12835 527 13010
rect 718 12835 781 13010
rect 2301 12911 2369 14827
rect 2828 12890 2884 15895
rect 3490 14970 3511 15755
rect 3511 14970 3553 15755
rect 3553 14970 3569 15755
rect 3490 14962 3569 14970
rect 15881 15505 15982 15917
rect 3332 12909 3400 14825
rect 12639 12660 12881 13073
rect -36 11330 95 12090
rect 197 10324 268 12084
rect 455 9380 526 11152
rect 713 10324 784 12084
rect 971 9380 1042 11152
rect 1229 10324 1300 12084
rect 1487 9380 1558 11152
rect 1745 10324 1816 12084
rect 2003 9380 2074 11152
rect 2261 10324 2332 12084
rect 2519 9380 2590 11152
rect 2777 10324 2848 12084
rect 3035 9380 3106 11152
rect 3293 10324 3364 12084
rect 3472 11329 3603 12089
rect 8065 9675 8155 9765
rect 8065 8985 8155 9075
rect 4886 4935 4966 5015
rect 6382 5125 6472 5215
rect -44 4495 76 4615
rect 3182 4495 3302 4615
rect 8070 5000 8150 5080
rect 15882 8978 15982 9078
rect 19896 5867 20144 6891
rect 15881 4701 15981 4801
rect 16760 5180 16860 5280
rect 19500 5180 19914 5280
rect -44 4260 76 4380
rect -297 2478 -256 3381
rect -256 2478 -190 3381
rect -190 2478 -21 3381
rect 3535 4275 3625 4365
rect 4474 302 4764 395
rect 6180 325 6317 377
rect 6717 4276 6807 4366
rect 9900 4270 9990 4360
rect 13080 4270 13170 4360
rect 15937 4270 16037 4370
rect 9358 495 9430 548
rect 7663 322 7955 374
rect 13604 20 13703 151
rect 6376 -139 6496 -27
rect 17213 322 17493 374
rect 18930 325 19040 377
rect 16101 -125 16181 -35
rect -80 -676 -20 -616
rect 3546 -3722 3626 -3642
rect -73 -3915 27 -3815
rect 880 -4945 980 -4845
rect 1524 -4944 1624 -4844
rect 2415 -4946 2515 -4846
rect 5987 -3723 6107 -3603
rect 3830 -4945 3930 -4845
rect 3547 -5212 3627 -5132
rect 16090 -3710 16190 -3610
rect 10022 -3915 10122 -3815
rect 16090 -4713 16190 -4613
rect 6273 -4946 6373 -4846
rect 10979 -4945 11079 -4845
rect 11621 -4946 11721 -4846
rect 12513 -4946 12613 -4846
rect 13928 -4946 14028 -4846
rect 16370 -4946 16470 -4846
rect 9845 -5205 9935 -5115
rect 10246 -5205 10336 -5115
rect 10245 -5613 10754 -5463
rect -90 -5755 -10 -5675
rect 62 -6580 267 -6500
rect 10970 -6573 11087 -6506
rect 62 -6720 267 -6640
rect 11612 -6713 11729 -6646
rect 62 -6860 267 -6780
rect 12504 -6854 12621 -6787
rect 62 -7000 267 -6920
rect 13920 -6993 14037 -6926
rect 62 -7140 267 -7060
rect 16363 -7134 16480 -7067
rect 880 -8805 980 -8705
rect -74 -8984 26 -8884
rect 1521 -8805 1621 -8705
rect 2415 -8805 2515 -8705
rect 3536 -8817 3636 -8717
rect 3832 -8819 3932 -8719
rect 6275 -8819 6375 -8719
rect 10022 -8983 10122 -8883
rect 3550 -9767 3620 -9697
rect 20101 -9760 20207 -9700
<< metal2 >>
rect -2716 17631 -2183 17909
rect -2023 17631 -1996 17909
rect -2718 17154 -2707 17433
rect -2559 17154 -1181 17433
rect -1033 17154 -1018 17433
rect -2751 16410 -2378 16466
rect -2244 16410 -2234 16466
rect 2401 16331 2736 16335
rect 2401 16322 2421 16331
rect -654 16266 2421 16322
rect -1691 14601 -1238 14618
rect -1691 14507 -1675 14601
rect -1260 14572 -1238 14601
rect -654 14572 -598 16266
rect 2401 16260 2421 16266
rect 2717 16260 2736 16331
rect 2401 16254 2736 16260
rect 2807 15895 2900 15911
rect 2807 15783 2828 15895
rect -323 14936 -313 15783
rect -134 15763 2828 15783
rect -134 14970 2131 15763
rect 2210 14970 2828 15763
rect -134 14936 2828 14970
rect -1260 14516 -598 14572
rect 2253 14827 2404 14859
rect -1260 14507 -1238 14516
rect -1691 14492 -1238 14507
rect -2751 13914 -2378 13970
rect -2244 13914 -2234 13970
rect 2253 13293 2301 14827
rect 177 13126 2301 13293
rect 177 13010 283 13126
rect 177 12835 197 13010
rect 260 12835 283 13010
rect 177 12819 283 12835
rect 393 13010 599 13023
rect 393 12835 464 13010
rect 527 12835 599 13010
rect -1691 12105 -1238 12122
rect 393 12107 599 12835
rect 698 13010 804 13126
rect 698 12835 718 13010
rect 781 12835 804 13010
rect 2253 12911 2301 13126
rect 2369 12911 2404 14827
rect 2253 12886 2404 12911
rect 2565 12890 2828 14936
rect 2884 15783 2900 15895
rect 2884 15755 3589 15783
rect 2884 14962 3490 15755
rect 3569 14962 3589 15755
rect 2884 14936 3589 14962
rect 2884 12890 3141 14936
rect 3319 14849 3412 14853
rect 2288 12882 2381 12886
rect 2565 12865 3141 12890
rect 3296 14847 3447 14849
rect 3754 14847 3945 20708
rect 19045 19437 19165 19448
rect 19045 19020 19052 19437
rect 19158 19020 19165 19437
rect 16605 16596 16865 16607
rect 16605 16176 16610 16596
rect 16859 16176 16865 16596
rect 3296 14825 3945 14847
rect 3296 12909 3332 14825
rect 3400 14656 3945 14825
rect 15872 15917 15992 15928
rect 15872 15505 15881 15917
rect 15982 15505 15992 15917
rect 3400 12909 3447 14656
rect 3296 12876 3447 12909
rect 12631 13073 12891 13084
rect 2807 12864 2900 12865
rect 698 12826 804 12835
rect 12631 12660 12639 13073
rect 12881 12660 12891 13073
rect -1691 12011 -1675 12105
rect -1260 12011 -1238 12105
rect -1691 11996 -1238 12011
rect -918 12090 3657 12107
rect -918 12089 -36 12090
rect -2751 11418 -2378 11474
rect -2244 11418 -2234 11474
rect -1350 10388 -1282 11996
rect -918 11332 -888 12089
rect -388 11332 -36 12089
rect -918 11330 -36 11332
rect 95 12089 3657 12090
rect 95 12084 3472 12089
rect 95 11330 197 12084
rect -918 11310 197 11330
rect -1350 10320 -574 10388
rect -1691 9609 -1238 9626
rect -1691 9515 -1675 9609
rect -1260 9580 -1238 9609
rect -1260 9524 -686 9580
rect -1260 9515 -1238 9524
rect -1691 9500 -1238 9515
rect -2751 8922 -2378 8978
rect -2244 8922 -2234 8978
rect -1691 7113 -1238 7130
rect -1691 7019 -1675 7113
rect -1260 7084 -1238 7113
rect -1260 7028 -798 7084
rect -1260 7019 -1238 7028
rect -1691 7004 -1238 7019
rect -1987 6896 -1744 6914
rect -2751 6426 -2378 6482
rect -2244 6426 -2234 6482
rect -1987 5851 -1971 6896
rect -1769 5851 -1744 6896
rect -1987 5826 -1744 5851
rect -1691 4617 -1238 4634
rect -1691 4523 -1675 4617
rect -1260 4588 -1238 4617
rect -1260 4532 -910 4588
rect -1260 4523 -1238 4532
rect -1691 4508 -1238 4523
rect -2751 3930 -2378 3986
rect -2244 3930 -2234 3986
rect -1691 2121 -1238 2138
rect -1691 2027 -1675 2121
rect -1260 2092 -1238 2121
rect -1260 2036 -1022 2092
rect -1260 2027 -1238 2036
rect -1691 2012 -1238 2027
rect -2751 1434 -2378 1490
rect -2244 1434 -2234 1490
rect -1691 -375 -1238 -358
rect -1691 -469 -1675 -375
rect -1260 -404 -1238 -375
rect -1260 -460 -1140 -404
rect -1260 -469 -1238 -460
rect -1691 -484 -1238 -469
rect -2751 -1062 -2378 -1006
rect -2244 -1062 -2234 -1006
rect -1691 -2871 -1257 -2854
rect -1691 -2965 -1675 -2871
rect -1260 -2965 -1257 -2871
rect -1691 -2980 -1257 -2965
rect -2751 -3558 -2378 -3502
rect -2244 -3558 -2234 -3502
rect -1313 -5247 -1257 -2980
rect -1196 -5083 -1140 -460
rect -1078 -4400 -1022 2036
rect -966 -4288 -910 4532
rect -854 -4184 -798 7028
rect -742 -4077 -686 9524
rect -630 -3958 -574 10320
rect 268 11310 713 12084
rect 197 10311 268 10324
rect 419 11152 541 11183
rect 419 9380 455 11152
rect 526 9380 541 11152
rect 784 11310 1229 12084
rect 713 10311 784 10324
rect 935 11152 1057 11183
rect 419 9302 541 9380
rect 935 9380 971 11152
rect 1042 9380 1057 11152
rect 1300 11310 1745 12084
rect 1229 10311 1300 10324
rect 1451 11152 1573 11183
rect 935 9302 1057 9380
rect 1451 9380 1487 11152
rect 1558 9380 1573 11152
rect 1816 11310 2261 12084
rect 1745 10311 1816 10324
rect 1967 11152 2089 11183
rect 1451 9302 1573 9380
rect 1967 9380 2003 11152
rect 2074 9380 2089 11152
rect 2332 11310 2777 12084
rect 2261 10311 2332 10324
rect 2483 11152 2605 11183
rect 1967 9302 2089 9380
rect 2483 9847 2519 11152
rect 2590 9847 2605 11152
rect 2848 11310 3293 12084
rect 2777 10311 2848 10324
rect 2999 11152 3121 11183
rect 2483 9321 2494 9847
rect 2594 9321 2605 9847
rect 2483 9302 2605 9321
rect 2999 10039 3035 11152
rect 3106 10039 3121 11152
rect 3364 11329 3472 12084
rect 3603 11329 3657 12089
rect 3364 11310 3657 11329
rect 3293 10311 3364 10324
rect 2999 9465 3009 10039
rect 3109 9465 3121 10039
rect 2999 9380 3035 9465
rect 3106 9380 3121 9465
rect 2999 9302 3121 9380
rect 8049 9765 8169 9780
rect 8049 9675 8065 9765
rect 8155 9675 8169 9765
rect 444 8672 515 9302
rect 957 8845 1028 9302
rect 1475 9061 1546 9302
rect 1995 9226 2066 9302
rect 1995 9155 7040 9226
rect 1475 8990 6770 9061
rect 957 8774 6510 8845
rect 444 8601 3298 8672
rect 3227 7637 3298 8601
rect 2737 7566 3298 7637
rect 2737 5663 2808 7566
rect 3227 7563 3298 7566
rect 6439 7362 6510 8774
rect 6699 8697 6770 8990
rect 6969 8883 7040 9155
rect 8049 9075 8169 9675
rect 8049 8985 8065 9075
rect 8155 8985 8169 9075
rect 8049 8970 8169 8985
rect 6969 8812 11293 8883
rect 6699 8626 9690 8697
rect 9619 7362 9690 8626
rect 11222 7772 11293 8812
rect 12631 8148 12891 12660
rect 14046 9335 14518 9346
rect 14046 9268 14069 9335
rect 14502 9268 14518 9335
rect 14046 9259 14518 9268
rect 11972 7888 12891 8148
rect 11222 7701 12034 7772
rect 11963 7362 12034 7701
rect 14447 7738 14518 9259
rect 15872 9078 15992 15505
rect 15872 8978 15882 9078
rect 15982 8978 15992 9078
rect 15872 8970 15992 8978
rect 16605 8959 16865 16176
rect 17140 9524 17659 9530
rect 17140 9458 17151 9524
rect 17642 9458 17659 9524
rect 17140 9453 17659 9458
rect 16605 8857 16864 8959
rect 15810 8597 16864 8857
rect 15810 8148 16070 8597
rect 15156 7888 16070 8148
rect 14447 7667 15620 7738
rect 17587 7721 17658 9453
rect 6439 7291 6746 7362
rect 9619 7291 9946 7362
rect 11963 7291 13126 7362
rect 1965 5592 2808 5663
rect -44 5121 76 5130
rect -44 4615 76 5001
rect 1965 4670 2036 5592
rect 3800 5220 6486 5230
rect 3800 5120 3810 5220
rect 3910 5215 6486 5220
rect 3910 5125 6382 5215
rect 6472 5125 6486 5215
rect 3910 5120 6486 5125
rect 3800 5110 6486 5120
rect 4875 5015 4979 5030
rect 4875 4935 4886 5015
rect 4966 4935 4979 5015
rect -50 4495 -44 4615
rect 76 4495 82 4615
rect 1965 4599 2291 4670
rect -44 4483 76 4495
rect -44 4380 76 4399
rect -44 3983 76 4260
rect -44 3854 76 3863
rect 2220 3464 2291 4599
rect 3165 4495 3182 4615
rect 3302 4495 3315 4615
rect 3165 4494 3310 4495
rect 4875 4372 4979 4935
rect 6675 4847 6746 7291
rect 3527 4365 4979 4372
rect 3527 4275 3535 4365
rect 3625 4275 4979 4365
rect 3527 4268 4979 4275
rect 6330 4776 6746 4847
rect 8058 5080 8160 5090
rect 8058 5000 8070 5080
rect 8150 5000 8160 5080
rect 2994 3780 3230 4043
rect 3067 3766 3230 3780
rect 3067 3603 3569 3766
rect -315 3381 4 3403
rect -315 2478 -297 3381
rect -21 2478 4 3381
rect -315 2453 4 2478
rect 3406 658 3569 3603
rect 6330 3564 6401 4776
rect 8058 4372 8160 5000
rect 9875 4847 9946 7291
rect 13055 4847 13126 7291
rect 6710 4366 8160 4372
rect 6710 4276 6717 4366
rect 6807 4276 8160 4366
rect 6710 4270 8160 4276
rect 9510 4776 9946 4847
rect 12690 4776 13126 4847
rect 9510 3564 9581 4776
rect 9890 4360 12183 4370
rect 9890 4270 9900 4360
rect 9990 4270 12183 4360
rect 9890 4260 12183 4270
rect 12690 3564 12761 4776
rect 13071 4360 15349 4370
rect 13071 4270 13080 4360
rect 13170 4270 15349 4360
rect 13071 4261 15349 4270
rect 15549 4198 15620 7667
rect 16521 7650 17658 7721
rect 15872 4801 15992 4810
rect 15872 4701 15881 4801
rect 15981 4701 15992 4801
rect 15872 4370 15992 4701
rect 16521 4664 16592 7650
rect 19045 7352 19165 19020
rect 18628 7232 19165 7352
rect 18628 5290 18748 7232
rect 19861 6891 20180 6914
rect 19861 5867 19896 6891
rect 20144 5867 20180 6891
rect 19861 5839 20180 5867
rect 16750 5280 19924 5290
rect 16750 5180 16760 5280
rect 16860 5180 19500 5280
rect 19914 5180 19924 5280
rect 16750 5170 19924 5180
rect 16521 4593 18199 4664
rect 15872 4270 15937 4370
rect 16037 4270 16046 4370
rect 15872 4261 16046 4270
rect 15872 4260 15992 4261
rect 15549 4127 15941 4198
rect 15870 3564 15941 4127
rect 6008 3493 6401 3564
rect 9188 3493 9581 3564
rect 12368 3493 12761 3564
rect 15548 3493 15941 3564
rect 18128 3478 18199 4593
rect 18586 3786 20575 4043
rect 3067 526 3569 658
rect 3067 243 3076 526
rect 3222 495 3569 526
rect 9285 548 9439 566
rect 9285 495 9358 548
rect 9430 495 9439 548
rect 3222 243 3231 495
rect 9285 454 9439 495
rect 4459 395 4880 409
rect 4459 302 4474 395
rect 4764 302 4880 395
rect 4459 291 4880 302
rect 3067 234 3231 243
rect 4764 285 4880 291
rect 6103 377 6333 387
rect 6103 325 6180 377
rect 6317 325 6333 377
rect 6103 285 6333 325
rect 4764 169 6333 285
rect 7644 374 8064 410
rect 7644 322 7663 374
rect 7955 322 8064 374
rect 7644 284 8064 322
rect 17195 374 17616 409
rect 17195 322 17213 374
rect 17493 322 17616 374
rect 17195 284 17616 322
rect 18839 377 19050 387
rect 18839 325 18930 377
rect 19040 325 19050 377
rect 18839 284 19050 325
rect 17195 231 19050 284
rect 4764 152 4844 169
rect 1561 72 4844 152
rect 9504 151 13713 163
rect 9504 106 13604 151
rect 1564 -607 1644 72
rect 9170 20 13604 106
rect 13703 20 13713 151
rect 17419 106 19050 231
rect 9170 10 13713 20
rect 3522 -139 6376 -27
rect 6496 -139 6506 -27
rect -451 -616 1644 -607
rect -451 -676 -80 -616
rect -20 -676 1644 -616
rect -451 -687 1644 -676
rect 3523 -3642 3645 -139
rect 9170 -227 9323 10
rect 3523 -3722 3546 -3642
rect 3626 -3722 3645 -3642
rect 3523 -3733 3645 -3722
rect 5970 -380 9323 -227
rect 16080 -35 16200 -26
rect 16080 -125 16101 -35
rect 16181 -125 16200 -35
rect 5970 -3603 6123 -380
rect 5970 -3723 5987 -3603
rect 6107 -3723 6123 -3603
rect 16080 -3610 16200 -125
rect 16080 -3710 16090 -3610
rect 16190 -3710 16200 -3610
rect 16080 -3720 16200 -3710
rect 5970 -3740 6123 -3723
rect -90 -3815 10136 -3800
rect -90 -3915 -73 -3815
rect 27 -3915 10022 -3815
rect 10122 -3915 10136 -3815
rect -90 -3930 10136 -3915
rect -635 -4038 140 -3958
rect -635 -4077 140 -4066
rect -742 -4133 140 -4077
rect -635 -4146 140 -4133
rect -635 -4184 140 -4174
rect -854 -4240 140 -4184
rect -635 -4254 140 -4240
rect -635 -4288 140 -4282
rect -966 -4344 140 -4288
rect -635 -4362 140 -4344
rect -635 -4400 140 -4390
rect -1078 -4456 140 -4400
rect -635 -4470 140 -4456
rect 16080 -4613 16200 -4606
rect 16080 -4713 16090 -4613
rect 16190 -4713 16200 -4613
rect 16080 -4720 16200 -4713
rect 866 -4845 996 -4830
rect 866 -4945 880 -4845
rect 980 -4945 996 -4845
rect -1196 -5139 -957 -5083
rect -1313 -5303 -1069 -5247
rect -1691 -5367 -1181 -5350
rect -1691 -5461 -1675 -5367
rect -1260 -5461 -1181 -5367
rect -1691 -5476 -1181 -5461
rect -2751 -6054 -2378 -5998
rect -2244 -6054 -2234 -5998
rect -1237 -6779 -1181 -5476
rect -1125 -6657 -1069 -5303
rect -1013 -6514 -957 -5139
rect -461 -5689 -90 -5675
rect -463 -5745 -90 -5689
rect -461 -5755 -90 -5745
rect -629 -6514 62 -6500
rect -1013 -6570 62 -6514
rect -629 -6580 62 -6570
rect 267 -6580 289 -6500
rect -629 -6657 62 -6640
rect -1125 -6713 62 -6657
rect -629 -6720 62 -6713
rect 267 -6720 289 -6640
rect -1237 -6780 -579 -6779
rect -1237 -6835 62 -6780
rect -629 -6860 62 -6835
rect 267 -6860 289 -6780
rect -629 -6940 62 -6920
rect -714 -6996 62 -6940
rect -1691 -7863 -1238 -7846
rect -1691 -7957 -1675 -7863
rect -1260 -7892 -1238 -7863
rect -714 -7892 -658 -6996
rect -629 -7000 62 -6996
rect 267 -7000 289 -6920
rect -629 -7140 62 -7060
rect 267 -7140 289 -7060
rect -1260 -7948 -658 -7892
rect -1260 -7957 -1238 -7948
rect -1691 -7972 -1238 -7957
rect -2751 -8550 -2378 -8494
rect -2244 -8550 -2234 -8494
rect -1691 -10359 -1238 -10342
rect -1691 -10453 -1675 -10359
rect -1260 -10388 -1238 -10359
rect -613 -10388 -557 -7140
rect 866 -8705 996 -4945
rect 866 -8805 880 -8705
rect 980 -8805 996 -8705
rect 866 -8820 996 -8805
rect 1508 -4844 1638 -4830
rect 1508 -4944 1524 -4844
rect 1624 -4944 1638 -4844
rect 1508 -8705 1638 -4944
rect 1508 -8805 1521 -8705
rect 1621 -8805 1638 -8705
rect 1508 -8820 1638 -8805
rect 2400 -4846 2530 -4830
rect 2400 -4946 2415 -4846
rect 2515 -4946 2530 -4846
rect 2400 -8705 2530 -4946
rect 3816 -4845 3946 -4830
rect 3816 -4945 3830 -4845
rect 3930 -4945 3946 -4845
rect 2400 -8805 2415 -8705
rect 2515 -8805 2530 -8705
rect 2400 -8820 2530 -8805
rect 3523 -5132 3646 -5117
rect 3523 -5212 3547 -5132
rect 3627 -5212 3646 -5132
rect 3523 -8717 3646 -5212
rect 3523 -8817 3536 -8717
rect 3636 -8817 3646 -8717
rect 3523 -8829 3646 -8817
rect 3816 -8719 3946 -4945
rect 3816 -8819 3832 -8719
rect 3932 -8819 3946 -8719
rect 3816 -8829 3946 -8819
rect 6259 -4846 6389 -4830
rect 6259 -4946 6273 -4846
rect 6373 -4946 6389 -4846
rect 6259 -8719 6389 -4946
rect 10963 -4845 11093 -4830
rect 10963 -4945 10979 -4845
rect 11079 -4945 11093 -4845
rect 9820 -5115 10363 -5092
rect 9820 -5205 9845 -5115
rect 9935 -5205 10246 -5115
rect 10336 -5205 10363 -5115
rect 9820 -5232 10363 -5205
rect 10224 -5463 10778 -5447
rect 10224 -5613 10245 -5463
rect 10754 -5613 10778 -5463
rect 10224 -5631 10778 -5613
rect 6259 -8819 6275 -8719
rect 6375 -8819 6389 -8719
rect 6259 -8829 6389 -8819
rect 10963 -6506 11093 -4945
rect 10963 -6573 10970 -6506
rect 11087 -6573 11093 -6506
rect -90 -8883 10136 -8868
rect -90 -8884 10022 -8883
rect -90 -8984 -74 -8884
rect 26 -8983 10022 -8884
rect 10122 -8983 10136 -8883
rect 26 -8984 10136 -8983
rect -90 -8998 10136 -8984
rect -90 -9106 140 -9026
rect 10963 -9106 11093 -6573
rect 11605 -4846 11735 -4830
rect 11605 -4946 11621 -4846
rect 11721 -4946 11735 -4846
rect 11605 -6646 11735 -4946
rect 11605 -6713 11612 -6646
rect 11729 -6713 11735 -6646
rect -90 -9214 140 -9134
rect 11605 -9214 11735 -6713
rect 12497 -4846 12627 -4830
rect 12497 -4946 12513 -4846
rect 12613 -4946 12627 -4846
rect 12497 -6787 12627 -4946
rect 12497 -6854 12504 -6787
rect 12621 -6854 12627 -6787
rect -90 -9322 140 -9242
rect 12497 -9322 12627 -6854
rect 13913 -4846 14043 -4830
rect 13913 -4946 13928 -4846
rect 14028 -4946 14043 -4846
rect 13913 -6926 14043 -4946
rect 13913 -6993 13920 -6926
rect 14037 -6993 14043 -6926
rect -90 -9430 140 -9350
rect 13913 -9430 14043 -6993
rect 16356 -4846 16486 -4830
rect 16356 -4946 16370 -4846
rect 16470 -4946 16486 -4846
rect 16356 -7067 16486 -4946
rect 16356 -7134 16363 -7067
rect 16480 -7134 16486 -7067
rect -90 -9538 140 -9458
rect 16356 -9538 16486 -7134
rect 3541 -9697 3631 -9684
rect 3541 -9767 3550 -9697
rect 3620 -9767 3631 -9697
rect 19612 -9700 20214 -9694
rect 19612 -9760 20101 -9700
rect 20207 -9760 20214 -9700
rect 19612 -9766 20214 -9760
rect 3541 -9774 3631 -9767
rect -1260 -10444 -557 -10388
rect -1260 -10453 -1238 -10444
rect -1691 -10468 -1238 -10453
<< via2 >>
rect -888 11332 -388 12089
rect -1971 5851 -1769 6896
rect 2494 9380 2519 9847
rect 2519 9380 2590 9847
rect 2590 9380 2594 9847
rect 2494 9321 2594 9380
rect 3009 9465 3035 10039
rect 3035 9465 3106 10039
rect 3106 9465 3109 10039
rect 14069 9268 14502 9335
rect 17151 9458 17642 9524
rect -44 5001 76 5121
rect 3810 5120 3910 5220
rect -44 3863 76 3983
rect 3200 4504 3300 4604
rect 2544 3813 2677 4102
rect -297 2478 -21 3381
rect 19896 5867 20144 6891
rect 3076 243 3222 526
rect 10245 -5613 10754 -5463
<< metal3 >>
rect -913 12089 -358 12141
rect -913 11332 -888 12089
rect -388 11332 -358 12089
rect -1987 6913 -1744 6914
rect -913 6913 -358 11332
rect 3000 10039 3120 10051
rect 2485 9847 2605 9862
rect 2485 9321 2494 9847
rect 2594 9341 2605 9847
rect 3000 9465 3009 10039
rect 3109 9531 3120 10039
rect 3109 9524 17664 9531
rect 3109 9465 17151 9524
rect 3000 9458 17151 9465
rect 17642 9458 17664 9524
rect 3000 9452 17664 9458
rect 3000 9451 3120 9452
rect 2594 9335 14508 9341
rect 2594 9321 14069 9335
rect 2485 9268 14069 9321
rect 14502 9268 14508 9335
rect 2485 9262 14508 9268
rect -2707 6896 3188 6913
rect -2707 5851 -1971 6896
rect -1769 5851 3188 6896
rect -2707 5840 3188 5851
rect 19099 6891 20589 6913
rect 19099 5867 19896 6891
rect 20144 5867 20589 6891
rect 19099 5840 20589 5867
rect -1987 5826 -1744 5840
rect 3787 5220 3920 5230
rect -77 5121 86 5131
rect -2745 5001 -44 5121
rect 76 5001 86 5121
rect 3787 5120 3810 5220
rect 3910 5120 3920 5220
rect 3787 5110 3920 5120
rect -2745 4986 86 5001
rect -77 4982 86 4986
rect -172 4615 159 4623
rect 3797 4615 3917 5110
rect -2738 4604 3917 4615
rect -2738 4504 3200 4604
rect 3300 4504 3917 4604
rect -2738 4495 3917 4504
rect -172 4486 159 4495
rect 3190 4494 3330 4495
rect 6337 4394 6483 4617
rect -2744 4248 6483 4394
rect 2536 4102 2684 4125
rect 2536 3993 2544 4102
rect -62 3983 2544 3993
rect -62 3863 -44 3983
rect 76 3863 2544 3983
rect -62 3850 2544 3863
rect 2536 3813 2544 3850
rect 2677 3813 2684 4102
rect 2536 3791 2684 3813
rect -2719 3381 3 3403
rect -2719 2478 -297 3381
rect -21 2478 3 3381
rect -2719 2454 3 2478
rect 19105 2454 20529 3403
rect -315 2453 3 2454
rect 3067 526 3231 535
rect 3067 243 3076 526
rect 3222 243 3231 526
rect 3067 234 3231 243
rect 3076 -5466 3224 234
rect 10224 -5463 10778 -5447
rect 10224 -5466 10245 -5463
rect 3076 -5613 10245 -5466
rect 10754 -5613 10778 -5463
rect 3076 -5614 10778 -5613
rect 10224 -5631 10778 -5614
use ia_opamp  ia_opamp_0
timestamp 1720298254
transform 1 0 -3812 0 1 -243
box 3810 247 7000 9177
use sky130_fd_pr__nfet_g5v0d10v5_EHZ5KL  sky130_fd_pr__nfet_g5v0d10v5_EHZ5KL_0 paramcells
timestamp 1720214482
transform 1 0 2851 0 1 14380
box -715 -1802 715 1802
use sky130_fd_pr__pfet_g5v0d10v5_6HDYS4  sky130_fd_pr__pfet_g5v0d10v5_6HDYS4_0 paramcells
timestamp 1720214482
transform 1 0 491 0 1 12923
box -487 -397 487 397
use sky130_fd_pr__pfet_g5v0d10v5_SKQKSC  sky130_fd_pr__pfet_g5v0d10v5_SKQKSC_0 paramcells
timestamp 1720214482
transform -1 0 1781 0 -1 10729
box -1777 -1797 1777 1797
use sky130_fd_sc_hvl__decap_4  sky130_fd_sc_hvl__decap_4_0 $PDKPATH/libs.ref/sky130_fd_sc_hvl/mag
array 0 10 -2496 0 0 940
timestamp 1715205430
transform 0 1 -2684 -1 0 -7909
box -66 -43 450 897
use sky130_fd_sc_hvl__diode_2  sky130_fd_sc_hvl__diode_2_0 $PDKPATH/libs.ref/sky130_fd_sc_hvl/mag
array 0 10 -2496 0 0 -940
timestamp 1715205430
transform 0 -1 -1056 -1 0 -8101
box -66 -43 258 897
use sky130_fd_sc_hvl__fill_2  sky130_fd_sc_hvl__fill_2_0 $PDKPATH/libs.ref/sky130_fd_sc_hvl/mag
array 0 10 -2496 0 0 -940
timestamp 1715205430
transform 0 -1 -1056 -1 0 -7909
box -66 -43 258 897
use sky130_fd_sc_hvl__lsbuflv2hv_1  sky130_fd_sc_hvl__lsbuflv2hv_1_0 $PDKPATH/libs.ref/sky130_fd_sc_hvl/mag
array 0 10 -2496 0 0 1714
timestamp 1715205430
transform 0 1 -2684 -1 0 -8293
box -66 -43 2178 1671
use RB_array_20  x1
timestamp 1718246682
transform 1 0 -1780 0 1 -5002
box 1690 -194 11784 4950
use RB_array_20  x2
timestamp 1718246682
transform 1 0 -1780 0 1 -10070
box 1690 -194 11784 4950
use RB_array_20  x3
timestamp 1718246682
transform 1 0 8317 0 1 -5002
box 1690 -194 11784 4950
use ia_opamp  x4
timestamp 1720298254
transform 1 0 -628 0 1 -243
box 3810 247 7000 9177
use ia_opamp  x5
timestamp 1720298254
transform 1 0 2556 0 1 -243
box 3810 247 7000 9177
use ia_opamp  x6
timestamp 1720298254
transform 1 0 12108 0 1 -243
box 3810 247 7000 9177
use RB_array_20  x7
timestamp 1718246682
transform 1 0 8317 0 1 -10070
box 1690 -194 11784 4950
use ia_opamp  x8
timestamp 1720298254
transform 1 0 5740 0 1 -243
box 3810 247 7000 9177
use ia_opamp  x9
timestamp 1720298254
transform 1 0 8924 0 1 -243
box 3810 247 7000 9177
use sky130_fd_pr__res_high_po_0p69_WX3C5M  XR1 paramcells
timestamp 1718246682
transform 1 0 11794 0 1 10788
box -7606 -1804 7606 1804
use sky130_fd_pr__res_high_po_0p69_WX3C5M  XR2
timestamp 1718246682
transform -1 0 11794 0 -1 17792
box -7606 -1804 7606 1804
use sky130_fd_pr__res_high_po_0p69_WX3C5M  XR4
timestamp 1718246682
transform 1 0 11794 0 1 14290
box -7606 -1804 7606 1804
<< labels >>
flabel metal2 20316 3786 20575 4043 0 FreeSans 2400 0 0 0 VOUT
port 18 nsew
flabel dnwell -90 -5196 10004 -52 0 FreeSans 8000 0 0 0 x1
flabel dnwell 10007 -5196 20101 -52 0 FreeSans 8000 0 0 0 x3
flabel metal2 -461 -5755 -381 -5675 0 FreeSans 1600 0 0 0 AVOUT2
port 17 nsew
flabel dnwell -90 -10264 10004 -5120 0 FreeSans 8000 0 0 0 x2
flabel dnwell 10007 -10264 20101 -5120 0 FreeSans 8000 0 0 0 x7
flabel metal2 -451 -687 -371 -607 0 FreeSans 1600 0 0 0 AVOUT1
port 16 nsew
flabel dnwell 3188 8984 18400 12592 0 FreeSans 8000 0 0 0 XR1
flabel dnwell 15918 4 19108 8934 0 FreeSans 8000 0 0 0 x6
flabel dnwell 12734 4 15924 8934 0 FreeSans 8000 0 0 0 x9
flabel dnwell 9550 4 12740 8934 0 FreeSans 8000 0 0 0 x8
flabel dnwell 6366 4 9556 8934 0 FreeSans 8000 0 0 0 x5
flabel dnwell 3182 4 6372 8934 0 FreeSans 8000 0 0 0 x4
flabel dnwell 3188 12486 18400 16069 0 FreeSans 8000 0 0 0 XR4
flabel dnwell 4245 16050 19365 19553 0 FreeSans 8000 0 0 0 XR2
flabel metal2 -2351 17280 -2351 17280 0 FreeSans 1600 0 0 0 DVSS
port 20 nsew
flabel metal2 -2385 17763 -2385 17763 0 FreeSans 1600 0 0 0 DVDD
port 19 nsew
flabel metal2 -590 -7140 -510 -7060 0 FreeSans 960 0 0 0 D93v3
flabel metal2 -590 -7000 -510 -6920 0 FreeSans 960 0 0 0 D83v3
flabel metal2 -590 -6860 -510 -6780 0 FreeSans 960 0 0 0 D73v3
flabel metal2 -590 -6720 -510 -6640 0 FreeSans 960 0 0 0 D63v3
flabel metal2 -590 -6580 -510 -6500 0 FreeSans 960 0 0 0 D53v3
flabel metal2 -590 -4470 -510 -4390 0 FreeSans 960 0 0 0 D43v3
flabel metal2 -590 -4362 -510 -4282 0 FreeSans 960 0 0 0 D33v3
flabel metal2 -590 -4254 -510 -4174 0 FreeSans 960 0 0 0 D23v3
flabel metal2 -590 -4146 -510 -4066 0 FreeSans 960 0 0 0 D13v3
flabel metal2 -590 -4038 -510 -3958 0 FreeSans 960 0 0 0 D03v3
flabel metal2 -2751 -8550 -2378 -8494 0 FreeSans 960 0 0 0 D9
port 21 nsew
flabel metal2 -2751 -6054 -2378 -5998 0 FreeSans 960 0 0 0 D8
port 22 nsew
flabel metal2 -2751 -3558 -2378 -3502 0 FreeSans 960 0 0 0 D7
port 23 nsew
flabel metal2 -2751 -1062 -2378 -1006 0 FreeSans 960 0 0 0 D6
port 24 nsew
flabel metal2 -2751 1434 -2378 1490 0 FreeSans 960 0 0 0 D5
port 25 nsew
flabel metal2 -2751 3930 -2378 3986 0 FreeSans 960 0 0 0 D4
port 26 nsew
flabel metal2 -2751 6426 -2378 6482 0 FreeSans 960 0 0 0 D3
port 27 nsew
flabel metal2 -2751 8922 -2378 8978 0 FreeSans 960 0 0 0 D2
port 28 nsew
flabel metal2 -2751 11418 -2378 11474 0 FreeSans 960 0 0 0 D1
port 29 nsew
flabel metal2 -2751 13914 -2378 13970 0 FreeSans 960 0 0 0 D0
port 30 nsew
flabel metal2 -2751 16410 -2378 16466 0 FreeSans 960 0 0 0 ena
port 31 nsew
flabel metal3 -2744 4248 -2081 4394 0 FreeSans 960 0 0 0 V2
port 32 nsew
flabel metal3 -2738 4495 -2081 4615 0 FreeSans 960 0 0 0 V1
port 33 nsew
flabel metal3 -2745 4986 -2085 5121 0 FreeSans 960 0 0 0 G
port 34 nsew
flabel metal3 20378 5840 20589 6913 0 FreeSans 2400 90 0 0 VDD
port 35 nsew
flabel metal3 -2719 2454 -2551 3403 0 FreeSans 2400 90 0 0 VSS
port 36 nsew
flabel metal2 3754 20305 3945 20708 0 FreeSans 1600 90 0 0 ibias
port 37 nsew
<< end >>
