magic
tech sky130A
magscale 1 2
timestamp 1717127688
<< pwell >>
rect -1990 -1804 1990 1804
<< psubdiff >>
rect -1954 1734 -1858 1768
rect 1858 1734 1954 1768
rect -1954 1672 -1920 1734
rect 1920 1672 1954 1734
rect -1954 -1734 -1920 -1672
rect 1920 -1734 1954 -1672
rect -1954 -1768 -1858 -1734
rect 1858 -1768 1954 -1734
<< psubdiffcont >>
rect -1858 1734 1858 1768
rect -1954 -1672 -1920 1672
rect 1920 -1672 1954 1672
rect -1858 -1768 1858 -1734
<< xpolycontact >>
rect -1824 1206 -1686 1638
rect -1824 -1638 -1686 -1206
rect -1590 1206 -1452 1638
rect -1590 -1638 -1452 -1206
rect -1356 1206 -1218 1638
rect -1356 -1638 -1218 -1206
rect -1122 1206 -984 1638
rect -1122 -1638 -984 -1206
rect -888 1206 -750 1638
rect -888 -1638 -750 -1206
rect -654 1206 -516 1638
rect -654 -1638 -516 -1206
rect -420 1206 -282 1638
rect -420 -1638 -282 -1206
rect -186 1206 -48 1638
rect -186 -1638 -48 -1206
rect 48 1206 186 1638
rect 48 -1638 186 -1206
rect 282 1206 420 1638
rect 282 -1638 420 -1206
rect 516 1206 654 1638
rect 516 -1638 654 -1206
rect 750 1206 888 1638
rect 750 -1638 888 -1206
rect 984 1206 1122 1638
rect 984 -1638 1122 -1206
rect 1218 1206 1356 1638
rect 1218 -1638 1356 -1206
rect 1452 1206 1590 1638
rect 1452 -1638 1590 -1206
rect 1686 1206 1824 1638
rect 1686 -1638 1824 -1206
<< ppolyres >>
rect -1824 -1206 -1686 1206
rect -1590 -1206 -1452 1206
rect -1356 -1206 -1218 1206
rect -1122 -1206 -984 1206
rect -888 -1206 -750 1206
rect -654 -1206 -516 1206
rect -420 -1206 -282 1206
rect -186 -1206 -48 1206
rect 48 -1206 186 1206
rect 282 -1206 420 1206
rect 516 -1206 654 1206
rect 750 -1206 888 1206
rect 984 -1206 1122 1206
rect 1218 -1206 1356 1206
rect 1452 -1206 1590 1206
rect 1686 -1206 1824 1206
<< locali >>
rect -1954 1734 -1858 1768
rect 1858 1734 1954 1768
rect -1954 1672 -1920 1734
rect 1920 1672 1954 1734
rect -1954 -1734 -1920 -1672
rect 1920 -1734 1954 -1672
rect -1954 -1768 -1858 -1734
rect 1858 -1768 1954 -1734
<< viali >>
rect -1808 1223 -1702 1620
rect -1574 1223 -1468 1620
rect -1340 1223 -1234 1620
rect -1106 1223 -1000 1620
rect -872 1223 -766 1620
rect -638 1223 -532 1620
rect -404 1223 -298 1620
rect -170 1223 -64 1620
rect 64 1223 170 1620
rect 298 1223 404 1620
rect 532 1223 638 1620
rect 766 1223 872 1620
rect 1000 1223 1106 1620
rect 1234 1223 1340 1620
rect 1468 1223 1574 1620
rect 1702 1223 1808 1620
rect -1808 -1620 -1702 -1223
rect -1574 -1620 -1468 -1223
rect -1340 -1620 -1234 -1223
rect -1106 -1620 -1000 -1223
rect -872 -1620 -766 -1223
rect -638 -1620 -532 -1223
rect -404 -1620 -298 -1223
rect -170 -1620 -64 -1223
rect 64 -1620 170 -1223
rect 298 -1620 404 -1223
rect 532 -1620 638 -1223
rect 766 -1620 872 -1223
rect 1000 -1620 1106 -1223
rect 1234 -1620 1340 -1223
rect 1468 -1620 1574 -1223
rect 1702 -1620 1808 -1223
<< metal1 >>
rect -1814 1620 -1696 1632
rect -1814 1223 -1808 1620
rect -1702 1223 -1696 1620
rect -1814 1211 -1696 1223
rect -1580 1620 -1462 1632
rect -1580 1223 -1574 1620
rect -1468 1223 -1462 1620
rect -1580 1211 -1462 1223
rect -1346 1620 -1228 1632
rect -1346 1223 -1340 1620
rect -1234 1223 -1228 1620
rect -1346 1211 -1228 1223
rect -1112 1620 -994 1632
rect -1112 1223 -1106 1620
rect -1000 1223 -994 1620
rect -1112 1211 -994 1223
rect -878 1620 -760 1632
rect -878 1223 -872 1620
rect -766 1223 -760 1620
rect -878 1211 -760 1223
rect -644 1620 -526 1632
rect -644 1223 -638 1620
rect -532 1223 -526 1620
rect -644 1211 -526 1223
rect -410 1620 -292 1632
rect -410 1223 -404 1620
rect -298 1223 -292 1620
rect -410 1211 -292 1223
rect -176 1620 -58 1632
rect -176 1223 -170 1620
rect -64 1223 -58 1620
rect -176 1211 -58 1223
rect 58 1620 176 1632
rect 58 1223 64 1620
rect 170 1223 176 1620
rect 58 1211 176 1223
rect 292 1620 410 1632
rect 292 1223 298 1620
rect 404 1223 410 1620
rect 292 1211 410 1223
rect 526 1620 644 1632
rect 526 1223 532 1620
rect 638 1223 644 1620
rect 526 1211 644 1223
rect 760 1620 878 1632
rect 760 1223 766 1620
rect 872 1223 878 1620
rect 760 1211 878 1223
rect 994 1620 1112 1632
rect 994 1223 1000 1620
rect 1106 1223 1112 1620
rect 994 1211 1112 1223
rect 1228 1620 1346 1632
rect 1228 1223 1234 1620
rect 1340 1223 1346 1620
rect 1228 1211 1346 1223
rect 1462 1620 1580 1632
rect 1462 1223 1468 1620
rect 1574 1223 1580 1620
rect 1462 1211 1580 1223
rect 1696 1620 1814 1632
rect 1696 1223 1702 1620
rect 1808 1223 1814 1620
rect 1696 1211 1814 1223
rect -1814 -1223 -1696 -1211
rect -1814 -1620 -1808 -1223
rect -1702 -1620 -1696 -1223
rect -1814 -1632 -1696 -1620
rect -1580 -1223 -1462 -1211
rect -1580 -1620 -1574 -1223
rect -1468 -1620 -1462 -1223
rect -1580 -1632 -1462 -1620
rect -1346 -1223 -1228 -1211
rect -1346 -1620 -1340 -1223
rect -1234 -1620 -1228 -1223
rect -1346 -1632 -1228 -1620
rect -1112 -1223 -994 -1211
rect -1112 -1620 -1106 -1223
rect -1000 -1620 -994 -1223
rect -1112 -1632 -994 -1620
rect -878 -1223 -760 -1211
rect -878 -1620 -872 -1223
rect -766 -1620 -760 -1223
rect -878 -1632 -760 -1620
rect -644 -1223 -526 -1211
rect -644 -1620 -638 -1223
rect -532 -1620 -526 -1223
rect -644 -1632 -526 -1620
rect -410 -1223 -292 -1211
rect -410 -1620 -404 -1223
rect -298 -1620 -292 -1223
rect -410 -1632 -292 -1620
rect -176 -1223 -58 -1211
rect -176 -1620 -170 -1223
rect -64 -1620 -58 -1223
rect -176 -1632 -58 -1620
rect 58 -1223 176 -1211
rect 58 -1620 64 -1223
rect 170 -1620 176 -1223
rect 58 -1632 176 -1620
rect 292 -1223 410 -1211
rect 292 -1620 298 -1223
rect 404 -1620 410 -1223
rect 292 -1632 410 -1620
rect 526 -1223 644 -1211
rect 526 -1620 532 -1223
rect 638 -1620 644 -1223
rect 526 -1632 644 -1620
rect 760 -1223 878 -1211
rect 760 -1620 766 -1223
rect 872 -1620 878 -1223
rect 760 -1632 878 -1620
rect 994 -1223 1112 -1211
rect 994 -1620 1000 -1223
rect 1106 -1620 1112 -1223
rect 994 -1632 1112 -1620
rect 1228 -1223 1346 -1211
rect 1228 -1620 1234 -1223
rect 1340 -1620 1346 -1223
rect 1228 -1632 1346 -1620
rect 1462 -1223 1580 -1211
rect 1462 -1620 1468 -1223
rect 1574 -1620 1580 -1223
rect 1462 -1632 1580 -1620
rect 1696 -1223 1814 -1211
rect 1696 -1620 1702 -1223
rect 1808 -1620 1814 -1223
rect 1696 -1632 1814 -1620
<< properties >>
string FIXED_BBOX -1937 -1751 1937 1751
string gencell sky130_fd_pr__res_high_po_0p69
string library sky130
string parameters w 0.69 l 12.22 m 1 nx 16 wmin 0.690 lmin 0.50 rho 319.8 val 6.228k dummy 0 dw 0.0 term 194.82 sterm 0.0 caplen 0 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_high_po_0p35  sky130_fd_pr__res_high_po_0p69 sky130_fd_pr__res_high_po_1p41  sky130_fd_pr__res_high_po_2p85 sky130_fd_pr__res_high_po_5p73} snake 0 full_metal 1 wmax 0.690 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
