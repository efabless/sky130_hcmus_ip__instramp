magic
tech sky130A
magscale 1 2
timestamp 1717127688
<< pwell >>
rect -7606 -1804 7606 1804
<< psubdiff >>
rect -7570 1734 -7474 1768
rect 7474 1734 7570 1768
rect -7570 1672 -7536 1734
rect 7536 1672 7570 1734
rect -7570 -1734 -7536 -1672
rect 7536 -1734 7570 -1672
rect -7570 -1768 -7474 -1734
rect 7474 -1768 7570 -1734
<< psubdiffcont >>
rect -7474 1734 7474 1768
rect -7570 -1672 -7536 1672
rect 7536 -1672 7570 1672
rect -7474 -1768 7474 -1734
<< xpolycontact >>
rect -7440 1206 -7302 1638
rect -7440 -1638 -7302 -1206
rect -7206 1206 -7068 1638
rect -7206 -1638 -7068 -1206
rect -6972 1206 -6834 1638
rect -6972 -1638 -6834 -1206
rect -6738 1206 -6600 1638
rect -6738 -1638 -6600 -1206
rect -6504 1206 -6366 1638
rect -6504 -1638 -6366 -1206
rect -6270 1206 -6132 1638
rect -6270 -1638 -6132 -1206
rect -6036 1206 -5898 1638
rect -6036 -1638 -5898 -1206
rect -5802 1206 -5664 1638
rect -5802 -1638 -5664 -1206
rect -5568 1206 -5430 1638
rect -5568 -1638 -5430 -1206
rect -5334 1206 -5196 1638
rect -5334 -1638 -5196 -1206
rect -5100 1206 -4962 1638
rect -5100 -1638 -4962 -1206
rect -4866 1206 -4728 1638
rect -4866 -1638 -4728 -1206
rect -4632 1206 -4494 1638
rect -4632 -1638 -4494 -1206
rect -4398 1206 -4260 1638
rect -4398 -1638 -4260 -1206
rect -4164 1206 -4026 1638
rect -4164 -1638 -4026 -1206
rect -3930 1206 -3792 1638
rect -3930 -1638 -3792 -1206
rect -3696 1206 -3558 1638
rect -3696 -1638 -3558 -1206
rect -3462 1206 -3324 1638
rect -3462 -1638 -3324 -1206
rect -3228 1206 -3090 1638
rect -3228 -1638 -3090 -1206
rect -2994 1206 -2856 1638
rect -2994 -1638 -2856 -1206
rect -2760 1206 -2622 1638
rect -2760 -1638 -2622 -1206
rect -2526 1206 -2388 1638
rect -2526 -1638 -2388 -1206
rect -2292 1206 -2154 1638
rect -2292 -1638 -2154 -1206
rect -2058 1206 -1920 1638
rect -2058 -1638 -1920 -1206
rect -1824 1206 -1686 1638
rect -1824 -1638 -1686 -1206
rect -1590 1206 -1452 1638
rect -1590 -1638 -1452 -1206
rect -1356 1206 -1218 1638
rect -1356 -1638 -1218 -1206
rect -1122 1206 -984 1638
rect -1122 -1638 -984 -1206
rect -888 1206 -750 1638
rect -888 -1638 -750 -1206
rect -654 1206 -516 1638
rect -654 -1638 -516 -1206
rect -420 1206 -282 1638
rect -420 -1638 -282 -1206
rect -186 1206 -48 1638
rect -186 -1638 -48 -1206
rect 48 1206 186 1638
rect 48 -1638 186 -1206
rect 282 1206 420 1638
rect 282 -1638 420 -1206
rect 516 1206 654 1638
rect 516 -1638 654 -1206
rect 750 1206 888 1638
rect 750 -1638 888 -1206
rect 984 1206 1122 1638
rect 984 -1638 1122 -1206
rect 1218 1206 1356 1638
rect 1218 -1638 1356 -1206
rect 1452 1206 1590 1638
rect 1452 -1638 1590 -1206
rect 1686 1206 1824 1638
rect 1686 -1638 1824 -1206
rect 1920 1206 2058 1638
rect 1920 -1638 2058 -1206
rect 2154 1206 2292 1638
rect 2154 -1638 2292 -1206
rect 2388 1206 2526 1638
rect 2388 -1638 2526 -1206
rect 2622 1206 2760 1638
rect 2622 -1638 2760 -1206
rect 2856 1206 2994 1638
rect 2856 -1638 2994 -1206
rect 3090 1206 3228 1638
rect 3090 -1638 3228 -1206
rect 3324 1206 3462 1638
rect 3324 -1638 3462 -1206
rect 3558 1206 3696 1638
rect 3558 -1638 3696 -1206
rect 3792 1206 3930 1638
rect 3792 -1638 3930 -1206
rect 4026 1206 4164 1638
rect 4026 -1638 4164 -1206
rect 4260 1206 4398 1638
rect 4260 -1638 4398 -1206
rect 4494 1206 4632 1638
rect 4494 -1638 4632 -1206
rect 4728 1206 4866 1638
rect 4728 -1638 4866 -1206
rect 4962 1206 5100 1638
rect 4962 -1638 5100 -1206
rect 5196 1206 5334 1638
rect 5196 -1638 5334 -1206
rect 5430 1206 5568 1638
rect 5430 -1638 5568 -1206
rect 5664 1206 5802 1638
rect 5664 -1638 5802 -1206
rect 5898 1206 6036 1638
rect 5898 -1638 6036 -1206
rect 6132 1206 6270 1638
rect 6132 -1638 6270 -1206
rect 6366 1206 6504 1638
rect 6366 -1638 6504 -1206
rect 6600 1206 6738 1638
rect 6600 -1638 6738 -1206
rect 6834 1206 6972 1638
rect 6834 -1638 6972 -1206
rect 7068 1206 7206 1638
rect 7068 -1638 7206 -1206
rect 7302 1206 7440 1638
rect 7302 -1638 7440 -1206
<< ppolyres >>
rect -7440 -1206 -7302 1206
rect -7206 -1206 -7068 1206
rect -6972 -1206 -6834 1206
rect -6738 -1206 -6600 1206
rect -6504 -1206 -6366 1206
rect -6270 -1206 -6132 1206
rect -6036 -1206 -5898 1206
rect -5802 -1206 -5664 1206
rect -5568 -1206 -5430 1206
rect -5334 -1206 -5196 1206
rect -5100 -1206 -4962 1206
rect -4866 -1206 -4728 1206
rect -4632 -1206 -4494 1206
rect -4398 -1206 -4260 1206
rect -4164 -1206 -4026 1206
rect -3930 -1206 -3792 1206
rect -3696 -1206 -3558 1206
rect -3462 -1206 -3324 1206
rect -3228 -1206 -3090 1206
rect -2994 -1206 -2856 1206
rect -2760 -1206 -2622 1206
rect -2526 -1206 -2388 1206
rect -2292 -1206 -2154 1206
rect -2058 -1206 -1920 1206
rect -1824 -1206 -1686 1206
rect -1590 -1206 -1452 1206
rect -1356 -1206 -1218 1206
rect -1122 -1206 -984 1206
rect -888 -1206 -750 1206
rect -654 -1206 -516 1206
rect -420 -1206 -282 1206
rect -186 -1206 -48 1206
rect 48 -1206 186 1206
rect 282 -1206 420 1206
rect 516 -1206 654 1206
rect 750 -1206 888 1206
rect 984 -1206 1122 1206
rect 1218 -1206 1356 1206
rect 1452 -1206 1590 1206
rect 1686 -1206 1824 1206
rect 1920 -1206 2058 1206
rect 2154 -1206 2292 1206
rect 2388 -1206 2526 1206
rect 2622 -1206 2760 1206
rect 2856 -1206 2994 1206
rect 3090 -1206 3228 1206
rect 3324 -1206 3462 1206
rect 3558 -1206 3696 1206
rect 3792 -1206 3930 1206
rect 4026 -1206 4164 1206
rect 4260 -1206 4398 1206
rect 4494 -1206 4632 1206
rect 4728 -1206 4866 1206
rect 4962 -1206 5100 1206
rect 5196 -1206 5334 1206
rect 5430 -1206 5568 1206
rect 5664 -1206 5802 1206
rect 5898 -1206 6036 1206
rect 6132 -1206 6270 1206
rect 6366 -1206 6504 1206
rect 6600 -1206 6738 1206
rect 6834 -1206 6972 1206
rect 7068 -1206 7206 1206
rect 7302 -1206 7440 1206
<< locali >>
rect -7570 1734 -7474 1768
rect 7474 1734 7570 1768
rect -7570 1672 -7536 1734
rect 7536 1672 7570 1734
rect -7570 -1734 -7536 -1672
rect 7536 -1734 7570 -1672
rect -7570 -1768 -7474 -1734
rect 7474 -1768 7570 -1734
<< viali >>
rect -7424 1223 -7318 1620
rect -7190 1223 -7084 1620
rect -6956 1223 -6850 1620
rect -6722 1223 -6616 1620
rect -6488 1223 -6382 1620
rect -6254 1223 -6148 1620
rect -6020 1223 -5914 1620
rect -5786 1223 -5680 1620
rect -5552 1223 -5446 1620
rect -5318 1223 -5212 1620
rect -5084 1223 -4978 1620
rect -4850 1223 -4744 1620
rect -4616 1223 -4510 1620
rect -4382 1223 -4276 1620
rect -4148 1223 -4042 1620
rect -3914 1223 -3808 1620
rect -3680 1223 -3574 1620
rect -3446 1223 -3340 1620
rect -3212 1223 -3106 1620
rect -2978 1223 -2872 1620
rect -2744 1223 -2638 1620
rect -2510 1223 -2404 1620
rect -2276 1223 -2170 1620
rect -2042 1223 -1936 1620
rect -1808 1223 -1702 1620
rect -1574 1223 -1468 1620
rect -1340 1223 -1234 1620
rect -1106 1223 -1000 1620
rect -872 1223 -766 1620
rect -638 1223 -532 1620
rect -404 1223 -298 1620
rect -170 1223 -64 1620
rect 64 1223 170 1620
rect 298 1223 404 1620
rect 532 1223 638 1620
rect 766 1223 872 1620
rect 1000 1223 1106 1620
rect 1234 1223 1340 1620
rect 1468 1223 1574 1620
rect 1702 1223 1808 1620
rect 1936 1223 2042 1620
rect 2170 1223 2276 1620
rect 2404 1223 2510 1620
rect 2638 1223 2744 1620
rect 2872 1223 2978 1620
rect 3106 1223 3212 1620
rect 3340 1223 3446 1620
rect 3574 1223 3680 1620
rect 3808 1223 3914 1620
rect 4042 1223 4148 1620
rect 4276 1223 4382 1620
rect 4510 1223 4616 1620
rect 4744 1223 4850 1620
rect 4978 1223 5084 1620
rect 5212 1223 5318 1620
rect 5446 1223 5552 1620
rect 5680 1223 5786 1620
rect 5914 1223 6020 1620
rect 6148 1223 6254 1620
rect 6382 1223 6488 1620
rect 6616 1223 6722 1620
rect 6850 1223 6956 1620
rect 7084 1223 7190 1620
rect 7318 1223 7424 1620
rect -7424 -1620 -7318 -1223
rect -7190 -1620 -7084 -1223
rect -6956 -1620 -6850 -1223
rect -6722 -1620 -6616 -1223
rect -6488 -1620 -6382 -1223
rect -6254 -1620 -6148 -1223
rect -6020 -1620 -5914 -1223
rect -5786 -1620 -5680 -1223
rect -5552 -1620 -5446 -1223
rect -5318 -1620 -5212 -1223
rect -5084 -1620 -4978 -1223
rect -4850 -1620 -4744 -1223
rect -4616 -1620 -4510 -1223
rect -4382 -1620 -4276 -1223
rect -4148 -1620 -4042 -1223
rect -3914 -1620 -3808 -1223
rect -3680 -1620 -3574 -1223
rect -3446 -1620 -3340 -1223
rect -3212 -1620 -3106 -1223
rect -2978 -1620 -2872 -1223
rect -2744 -1620 -2638 -1223
rect -2510 -1620 -2404 -1223
rect -2276 -1620 -2170 -1223
rect -2042 -1620 -1936 -1223
rect -1808 -1620 -1702 -1223
rect -1574 -1620 -1468 -1223
rect -1340 -1620 -1234 -1223
rect -1106 -1620 -1000 -1223
rect -872 -1620 -766 -1223
rect -638 -1620 -532 -1223
rect -404 -1620 -298 -1223
rect -170 -1620 -64 -1223
rect 64 -1620 170 -1223
rect 298 -1620 404 -1223
rect 532 -1620 638 -1223
rect 766 -1620 872 -1223
rect 1000 -1620 1106 -1223
rect 1234 -1620 1340 -1223
rect 1468 -1620 1574 -1223
rect 1702 -1620 1808 -1223
rect 1936 -1620 2042 -1223
rect 2170 -1620 2276 -1223
rect 2404 -1620 2510 -1223
rect 2638 -1620 2744 -1223
rect 2872 -1620 2978 -1223
rect 3106 -1620 3212 -1223
rect 3340 -1620 3446 -1223
rect 3574 -1620 3680 -1223
rect 3808 -1620 3914 -1223
rect 4042 -1620 4148 -1223
rect 4276 -1620 4382 -1223
rect 4510 -1620 4616 -1223
rect 4744 -1620 4850 -1223
rect 4978 -1620 5084 -1223
rect 5212 -1620 5318 -1223
rect 5446 -1620 5552 -1223
rect 5680 -1620 5786 -1223
rect 5914 -1620 6020 -1223
rect 6148 -1620 6254 -1223
rect 6382 -1620 6488 -1223
rect 6616 -1620 6722 -1223
rect 6850 -1620 6956 -1223
rect 7084 -1620 7190 -1223
rect 7318 -1620 7424 -1223
<< metal1 >>
rect -7430 1620 -7312 1632
rect -7430 1223 -7424 1620
rect -7318 1223 -7312 1620
rect -7430 1211 -7312 1223
rect -7196 1620 -7078 1632
rect -7196 1223 -7190 1620
rect -7084 1223 -7078 1620
rect -7196 1211 -7078 1223
rect -6962 1620 -6844 1632
rect -6962 1223 -6956 1620
rect -6850 1223 -6844 1620
rect -6962 1211 -6844 1223
rect -6728 1620 -6610 1632
rect -6728 1223 -6722 1620
rect -6616 1223 -6610 1620
rect -6728 1211 -6610 1223
rect -6494 1620 -6376 1632
rect -6494 1223 -6488 1620
rect -6382 1223 -6376 1620
rect -6494 1211 -6376 1223
rect -6260 1620 -6142 1632
rect -6260 1223 -6254 1620
rect -6148 1223 -6142 1620
rect -6260 1211 -6142 1223
rect -6026 1620 -5908 1632
rect -6026 1223 -6020 1620
rect -5914 1223 -5908 1620
rect -6026 1211 -5908 1223
rect -5792 1620 -5674 1632
rect -5792 1223 -5786 1620
rect -5680 1223 -5674 1620
rect -5792 1211 -5674 1223
rect -5558 1620 -5440 1632
rect -5558 1223 -5552 1620
rect -5446 1223 -5440 1620
rect -5558 1211 -5440 1223
rect -5324 1620 -5206 1632
rect -5324 1223 -5318 1620
rect -5212 1223 -5206 1620
rect -5324 1211 -5206 1223
rect -5090 1620 -4972 1632
rect -5090 1223 -5084 1620
rect -4978 1223 -4972 1620
rect -5090 1211 -4972 1223
rect -4856 1620 -4738 1632
rect -4856 1223 -4850 1620
rect -4744 1223 -4738 1620
rect -4856 1211 -4738 1223
rect -4622 1620 -4504 1632
rect -4622 1223 -4616 1620
rect -4510 1223 -4504 1620
rect -4622 1211 -4504 1223
rect -4388 1620 -4270 1632
rect -4388 1223 -4382 1620
rect -4276 1223 -4270 1620
rect -4388 1211 -4270 1223
rect -4154 1620 -4036 1632
rect -4154 1223 -4148 1620
rect -4042 1223 -4036 1620
rect -4154 1211 -4036 1223
rect -3920 1620 -3802 1632
rect -3920 1223 -3914 1620
rect -3808 1223 -3802 1620
rect -3920 1211 -3802 1223
rect -3686 1620 -3568 1632
rect -3686 1223 -3680 1620
rect -3574 1223 -3568 1620
rect -3686 1211 -3568 1223
rect -3452 1620 -3334 1632
rect -3452 1223 -3446 1620
rect -3340 1223 -3334 1620
rect -3452 1211 -3334 1223
rect -3218 1620 -3100 1632
rect -3218 1223 -3212 1620
rect -3106 1223 -3100 1620
rect -3218 1211 -3100 1223
rect -2984 1620 -2866 1632
rect -2984 1223 -2978 1620
rect -2872 1223 -2866 1620
rect -2984 1211 -2866 1223
rect -2750 1620 -2632 1632
rect -2750 1223 -2744 1620
rect -2638 1223 -2632 1620
rect -2750 1211 -2632 1223
rect -2516 1620 -2398 1632
rect -2516 1223 -2510 1620
rect -2404 1223 -2398 1620
rect -2516 1211 -2398 1223
rect -2282 1620 -2164 1632
rect -2282 1223 -2276 1620
rect -2170 1223 -2164 1620
rect -2282 1211 -2164 1223
rect -2048 1620 -1930 1632
rect -2048 1223 -2042 1620
rect -1936 1223 -1930 1620
rect -2048 1211 -1930 1223
rect -1814 1620 -1696 1632
rect -1814 1223 -1808 1620
rect -1702 1223 -1696 1620
rect -1814 1211 -1696 1223
rect -1580 1620 -1462 1632
rect -1580 1223 -1574 1620
rect -1468 1223 -1462 1620
rect -1580 1211 -1462 1223
rect -1346 1620 -1228 1632
rect -1346 1223 -1340 1620
rect -1234 1223 -1228 1620
rect -1346 1211 -1228 1223
rect -1112 1620 -994 1632
rect -1112 1223 -1106 1620
rect -1000 1223 -994 1620
rect -1112 1211 -994 1223
rect -878 1620 -760 1632
rect -878 1223 -872 1620
rect -766 1223 -760 1620
rect -878 1211 -760 1223
rect -644 1620 -526 1632
rect -644 1223 -638 1620
rect -532 1223 -526 1620
rect -644 1211 -526 1223
rect -410 1620 -292 1632
rect -410 1223 -404 1620
rect -298 1223 -292 1620
rect -410 1211 -292 1223
rect -176 1620 -58 1632
rect -176 1223 -170 1620
rect -64 1223 -58 1620
rect -176 1211 -58 1223
rect 58 1620 176 1632
rect 58 1223 64 1620
rect 170 1223 176 1620
rect 58 1211 176 1223
rect 292 1620 410 1632
rect 292 1223 298 1620
rect 404 1223 410 1620
rect 292 1211 410 1223
rect 526 1620 644 1632
rect 526 1223 532 1620
rect 638 1223 644 1620
rect 526 1211 644 1223
rect 760 1620 878 1632
rect 760 1223 766 1620
rect 872 1223 878 1620
rect 760 1211 878 1223
rect 994 1620 1112 1632
rect 994 1223 1000 1620
rect 1106 1223 1112 1620
rect 994 1211 1112 1223
rect 1228 1620 1346 1632
rect 1228 1223 1234 1620
rect 1340 1223 1346 1620
rect 1228 1211 1346 1223
rect 1462 1620 1580 1632
rect 1462 1223 1468 1620
rect 1574 1223 1580 1620
rect 1462 1211 1580 1223
rect 1696 1620 1814 1632
rect 1696 1223 1702 1620
rect 1808 1223 1814 1620
rect 1696 1211 1814 1223
rect 1930 1620 2048 1632
rect 1930 1223 1936 1620
rect 2042 1223 2048 1620
rect 1930 1211 2048 1223
rect 2164 1620 2282 1632
rect 2164 1223 2170 1620
rect 2276 1223 2282 1620
rect 2164 1211 2282 1223
rect 2398 1620 2516 1632
rect 2398 1223 2404 1620
rect 2510 1223 2516 1620
rect 2398 1211 2516 1223
rect 2632 1620 2750 1632
rect 2632 1223 2638 1620
rect 2744 1223 2750 1620
rect 2632 1211 2750 1223
rect 2866 1620 2984 1632
rect 2866 1223 2872 1620
rect 2978 1223 2984 1620
rect 2866 1211 2984 1223
rect 3100 1620 3218 1632
rect 3100 1223 3106 1620
rect 3212 1223 3218 1620
rect 3100 1211 3218 1223
rect 3334 1620 3452 1632
rect 3334 1223 3340 1620
rect 3446 1223 3452 1620
rect 3334 1211 3452 1223
rect 3568 1620 3686 1632
rect 3568 1223 3574 1620
rect 3680 1223 3686 1620
rect 3568 1211 3686 1223
rect 3802 1620 3920 1632
rect 3802 1223 3808 1620
rect 3914 1223 3920 1620
rect 3802 1211 3920 1223
rect 4036 1620 4154 1632
rect 4036 1223 4042 1620
rect 4148 1223 4154 1620
rect 4036 1211 4154 1223
rect 4270 1620 4388 1632
rect 4270 1223 4276 1620
rect 4382 1223 4388 1620
rect 4270 1211 4388 1223
rect 4504 1620 4622 1632
rect 4504 1223 4510 1620
rect 4616 1223 4622 1620
rect 4504 1211 4622 1223
rect 4738 1620 4856 1632
rect 4738 1223 4744 1620
rect 4850 1223 4856 1620
rect 4738 1211 4856 1223
rect 4972 1620 5090 1632
rect 4972 1223 4978 1620
rect 5084 1223 5090 1620
rect 4972 1211 5090 1223
rect 5206 1620 5324 1632
rect 5206 1223 5212 1620
rect 5318 1223 5324 1620
rect 5206 1211 5324 1223
rect 5440 1620 5558 1632
rect 5440 1223 5446 1620
rect 5552 1223 5558 1620
rect 5440 1211 5558 1223
rect 5674 1620 5792 1632
rect 5674 1223 5680 1620
rect 5786 1223 5792 1620
rect 5674 1211 5792 1223
rect 5908 1620 6026 1632
rect 5908 1223 5914 1620
rect 6020 1223 6026 1620
rect 5908 1211 6026 1223
rect 6142 1620 6260 1632
rect 6142 1223 6148 1620
rect 6254 1223 6260 1620
rect 6142 1211 6260 1223
rect 6376 1620 6494 1632
rect 6376 1223 6382 1620
rect 6488 1223 6494 1620
rect 6376 1211 6494 1223
rect 6610 1620 6728 1632
rect 6610 1223 6616 1620
rect 6722 1223 6728 1620
rect 6610 1211 6728 1223
rect 6844 1620 6962 1632
rect 6844 1223 6850 1620
rect 6956 1223 6962 1620
rect 6844 1211 6962 1223
rect 7078 1620 7196 1632
rect 7078 1223 7084 1620
rect 7190 1223 7196 1620
rect 7078 1211 7196 1223
rect 7312 1620 7430 1632
rect 7312 1223 7318 1620
rect 7424 1223 7430 1620
rect 7312 1211 7430 1223
rect -7430 -1223 -7312 -1211
rect -7430 -1620 -7424 -1223
rect -7318 -1620 -7312 -1223
rect -7430 -1632 -7312 -1620
rect -7196 -1223 -7078 -1211
rect -7196 -1620 -7190 -1223
rect -7084 -1620 -7078 -1223
rect -7196 -1632 -7078 -1620
rect -6962 -1223 -6844 -1211
rect -6962 -1620 -6956 -1223
rect -6850 -1620 -6844 -1223
rect -6962 -1632 -6844 -1620
rect -6728 -1223 -6610 -1211
rect -6728 -1620 -6722 -1223
rect -6616 -1620 -6610 -1223
rect -6728 -1632 -6610 -1620
rect -6494 -1223 -6376 -1211
rect -6494 -1620 -6488 -1223
rect -6382 -1620 -6376 -1223
rect -6494 -1632 -6376 -1620
rect -6260 -1223 -6142 -1211
rect -6260 -1620 -6254 -1223
rect -6148 -1620 -6142 -1223
rect -6260 -1632 -6142 -1620
rect -6026 -1223 -5908 -1211
rect -6026 -1620 -6020 -1223
rect -5914 -1620 -5908 -1223
rect -6026 -1632 -5908 -1620
rect -5792 -1223 -5674 -1211
rect -5792 -1620 -5786 -1223
rect -5680 -1620 -5674 -1223
rect -5792 -1632 -5674 -1620
rect -5558 -1223 -5440 -1211
rect -5558 -1620 -5552 -1223
rect -5446 -1620 -5440 -1223
rect -5558 -1632 -5440 -1620
rect -5324 -1223 -5206 -1211
rect -5324 -1620 -5318 -1223
rect -5212 -1620 -5206 -1223
rect -5324 -1632 -5206 -1620
rect -5090 -1223 -4972 -1211
rect -5090 -1620 -5084 -1223
rect -4978 -1620 -4972 -1223
rect -5090 -1632 -4972 -1620
rect -4856 -1223 -4738 -1211
rect -4856 -1620 -4850 -1223
rect -4744 -1620 -4738 -1223
rect -4856 -1632 -4738 -1620
rect -4622 -1223 -4504 -1211
rect -4622 -1620 -4616 -1223
rect -4510 -1620 -4504 -1223
rect -4622 -1632 -4504 -1620
rect -4388 -1223 -4270 -1211
rect -4388 -1620 -4382 -1223
rect -4276 -1620 -4270 -1223
rect -4388 -1632 -4270 -1620
rect -4154 -1223 -4036 -1211
rect -4154 -1620 -4148 -1223
rect -4042 -1620 -4036 -1223
rect -4154 -1632 -4036 -1620
rect -3920 -1223 -3802 -1211
rect -3920 -1620 -3914 -1223
rect -3808 -1620 -3802 -1223
rect -3920 -1632 -3802 -1620
rect -3686 -1223 -3568 -1211
rect -3686 -1620 -3680 -1223
rect -3574 -1620 -3568 -1223
rect -3686 -1632 -3568 -1620
rect -3452 -1223 -3334 -1211
rect -3452 -1620 -3446 -1223
rect -3340 -1620 -3334 -1223
rect -3452 -1632 -3334 -1620
rect -3218 -1223 -3100 -1211
rect -3218 -1620 -3212 -1223
rect -3106 -1620 -3100 -1223
rect -3218 -1632 -3100 -1620
rect -2984 -1223 -2866 -1211
rect -2984 -1620 -2978 -1223
rect -2872 -1620 -2866 -1223
rect -2984 -1632 -2866 -1620
rect -2750 -1223 -2632 -1211
rect -2750 -1620 -2744 -1223
rect -2638 -1620 -2632 -1223
rect -2750 -1632 -2632 -1620
rect -2516 -1223 -2398 -1211
rect -2516 -1620 -2510 -1223
rect -2404 -1620 -2398 -1223
rect -2516 -1632 -2398 -1620
rect -2282 -1223 -2164 -1211
rect -2282 -1620 -2276 -1223
rect -2170 -1620 -2164 -1223
rect -2282 -1632 -2164 -1620
rect -2048 -1223 -1930 -1211
rect -2048 -1620 -2042 -1223
rect -1936 -1620 -1930 -1223
rect -2048 -1632 -1930 -1620
rect -1814 -1223 -1696 -1211
rect -1814 -1620 -1808 -1223
rect -1702 -1620 -1696 -1223
rect -1814 -1632 -1696 -1620
rect -1580 -1223 -1462 -1211
rect -1580 -1620 -1574 -1223
rect -1468 -1620 -1462 -1223
rect -1580 -1632 -1462 -1620
rect -1346 -1223 -1228 -1211
rect -1346 -1620 -1340 -1223
rect -1234 -1620 -1228 -1223
rect -1346 -1632 -1228 -1620
rect -1112 -1223 -994 -1211
rect -1112 -1620 -1106 -1223
rect -1000 -1620 -994 -1223
rect -1112 -1632 -994 -1620
rect -878 -1223 -760 -1211
rect -878 -1620 -872 -1223
rect -766 -1620 -760 -1223
rect -878 -1632 -760 -1620
rect -644 -1223 -526 -1211
rect -644 -1620 -638 -1223
rect -532 -1620 -526 -1223
rect -644 -1632 -526 -1620
rect -410 -1223 -292 -1211
rect -410 -1620 -404 -1223
rect -298 -1620 -292 -1223
rect -410 -1632 -292 -1620
rect -176 -1223 -58 -1211
rect -176 -1620 -170 -1223
rect -64 -1620 -58 -1223
rect -176 -1632 -58 -1620
rect 58 -1223 176 -1211
rect 58 -1620 64 -1223
rect 170 -1620 176 -1223
rect 58 -1632 176 -1620
rect 292 -1223 410 -1211
rect 292 -1620 298 -1223
rect 404 -1620 410 -1223
rect 292 -1632 410 -1620
rect 526 -1223 644 -1211
rect 526 -1620 532 -1223
rect 638 -1620 644 -1223
rect 526 -1632 644 -1620
rect 760 -1223 878 -1211
rect 760 -1620 766 -1223
rect 872 -1620 878 -1223
rect 760 -1632 878 -1620
rect 994 -1223 1112 -1211
rect 994 -1620 1000 -1223
rect 1106 -1620 1112 -1223
rect 994 -1632 1112 -1620
rect 1228 -1223 1346 -1211
rect 1228 -1620 1234 -1223
rect 1340 -1620 1346 -1223
rect 1228 -1632 1346 -1620
rect 1462 -1223 1580 -1211
rect 1462 -1620 1468 -1223
rect 1574 -1620 1580 -1223
rect 1462 -1632 1580 -1620
rect 1696 -1223 1814 -1211
rect 1696 -1620 1702 -1223
rect 1808 -1620 1814 -1223
rect 1696 -1632 1814 -1620
rect 1930 -1223 2048 -1211
rect 1930 -1620 1936 -1223
rect 2042 -1620 2048 -1223
rect 1930 -1632 2048 -1620
rect 2164 -1223 2282 -1211
rect 2164 -1620 2170 -1223
rect 2276 -1620 2282 -1223
rect 2164 -1632 2282 -1620
rect 2398 -1223 2516 -1211
rect 2398 -1620 2404 -1223
rect 2510 -1620 2516 -1223
rect 2398 -1632 2516 -1620
rect 2632 -1223 2750 -1211
rect 2632 -1620 2638 -1223
rect 2744 -1620 2750 -1223
rect 2632 -1632 2750 -1620
rect 2866 -1223 2984 -1211
rect 2866 -1620 2872 -1223
rect 2978 -1620 2984 -1223
rect 2866 -1632 2984 -1620
rect 3100 -1223 3218 -1211
rect 3100 -1620 3106 -1223
rect 3212 -1620 3218 -1223
rect 3100 -1632 3218 -1620
rect 3334 -1223 3452 -1211
rect 3334 -1620 3340 -1223
rect 3446 -1620 3452 -1223
rect 3334 -1632 3452 -1620
rect 3568 -1223 3686 -1211
rect 3568 -1620 3574 -1223
rect 3680 -1620 3686 -1223
rect 3568 -1632 3686 -1620
rect 3802 -1223 3920 -1211
rect 3802 -1620 3808 -1223
rect 3914 -1620 3920 -1223
rect 3802 -1632 3920 -1620
rect 4036 -1223 4154 -1211
rect 4036 -1620 4042 -1223
rect 4148 -1620 4154 -1223
rect 4036 -1632 4154 -1620
rect 4270 -1223 4388 -1211
rect 4270 -1620 4276 -1223
rect 4382 -1620 4388 -1223
rect 4270 -1632 4388 -1620
rect 4504 -1223 4622 -1211
rect 4504 -1620 4510 -1223
rect 4616 -1620 4622 -1223
rect 4504 -1632 4622 -1620
rect 4738 -1223 4856 -1211
rect 4738 -1620 4744 -1223
rect 4850 -1620 4856 -1223
rect 4738 -1632 4856 -1620
rect 4972 -1223 5090 -1211
rect 4972 -1620 4978 -1223
rect 5084 -1620 5090 -1223
rect 4972 -1632 5090 -1620
rect 5206 -1223 5324 -1211
rect 5206 -1620 5212 -1223
rect 5318 -1620 5324 -1223
rect 5206 -1632 5324 -1620
rect 5440 -1223 5558 -1211
rect 5440 -1620 5446 -1223
rect 5552 -1620 5558 -1223
rect 5440 -1632 5558 -1620
rect 5674 -1223 5792 -1211
rect 5674 -1620 5680 -1223
rect 5786 -1620 5792 -1223
rect 5674 -1632 5792 -1620
rect 5908 -1223 6026 -1211
rect 5908 -1620 5914 -1223
rect 6020 -1620 6026 -1223
rect 5908 -1632 6026 -1620
rect 6142 -1223 6260 -1211
rect 6142 -1620 6148 -1223
rect 6254 -1620 6260 -1223
rect 6142 -1632 6260 -1620
rect 6376 -1223 6494 -1211
rect 6376 -1620 6382 -1223
rect 6488 -1620 6494 -1223
rect 6376 -1632 6494 -1620
rect 6610 -1223 6728 -1211
rect 6610 -1620 6616 -1223
rect 6722 -1620 6728 -1223
rect 6610 -1632 6728 -1620
rect 6844 -1223 6962 -1211
rect 6844 -1620 6850 -1223
rect 6956 -1620 6962 -1223
rect 6844 -1632 6962 -1620
rect 7078 -1223 7196 -1211
rect 7078 -1620 7084 -1223
rect 7190 -1620 7196 -1223
rect 7078 -1632 7196 -1620
rect 7312 -1223 7430 -1211
rect 7312 -1620 7318 -1223
rect 7424 -1620 7430 -1223
rect 7312 -1632 7430 -1620
<< properties >>
string FIXED_BBOX -7553 -1751 7553 1751
string gencell sky130_fd_pr__res_high_po_0p69
string library sky130
string parameters w 0.69 l 12.22 m 1 nx 64 wmin 0.690 lmin 0.50 rho 319.8 val 6.228k dummy 0 dw 0.0 term 194.82 sterm 0.0 caplen 0 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_high_po_0p35  sky130_fd_pr__res_high_po_0p69 sky130_fd_pr__res_high_po_1p41  sky130_fd_pr__res_high_po_2p85 sky130_fd_pr__res_high_po_5p73} snake 0 full_metal 1 wmax 0.690 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
