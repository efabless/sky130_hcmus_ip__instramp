magic
tech sky130A
magscale 1 2
timestamp 1718246682
<< pwell >>
rect -235 -1804 235 1804
<< psubdiff >>
rect -199 1734 -103 1768
rect 103 1734 199 1768
rect -199 1672 -165 1734
rect 165 1672 199 1734
rect -199 -1734 -165 -1672
rect 165 -1734 199 -1672
rect -199 -1768 -103 -1734
rect 103 -1768 199 -1734
<< psubdiffcont >>
rect -103 1734 103 1768
rect -199 -1672 -165 1672
rect 165 -1672 199 1672
rect -103 -1768 103 -1734
<< xpolycontact >>
rect -69 1206 69 1638
rect -69 -1638 69 -1206
<< ppolyres >>
rect -69 -1206 69 1206
<< locali >>
rect -199 1734 -103 1768
rect 103 1734 199 1768
rect -199 1672 -165 1734
rect 165 1672 199 1734
rect -199 -1734 -165 -1672
rect 165 -1734 199 -1672
rect -199 -1768 -103 -1734
rect 103 -1768 199 -1734
<< viali >>
rect -53 1223 53 1620
rect -53 -1620 53 -1223
<< metal1 >>
rect -59 1620 59 1632
rect -59 1223 -53 1620
rect 53 1223 59 1620
rect -59 1211 59 1223
rect -59 -1223 59 -1211
rect -59 -1620 -53 -1223
rect 53 -1620 59 -1223
rect -59 -1632 59 -1620
<< properties >>
string FIXED_BBOX -182 -1751 182 1751
string gencell sky130_fd_pr__res_high_po_0p69
string library sky130
string parameters w 0.690 l 12.22 m 1 nx 1 wmin 0.690 lmin 0.50 rho 319.8 val 6.228k dummy 0 dw 0.0 term 194.82 sterm 0.0 caplen 0 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_high_po_0p35  sky130_fd_pr__res_high_po_0p69 sky130_fd_pr__res_high_po_1p41  sky130_fd_pr__res_high_po_2p85 sky130_fd_pr__res_high_po_5p73} snake 0 full_metal 1 wmax 0.690 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
