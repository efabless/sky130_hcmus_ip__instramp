magic
tech sky130A
magscale 1 2
timestamp 1716807968
<< pwell >>
rect -715 -1069 715 1069
<< mvnmos >>
rect -487 661 -287 811
rect -229 661 -29 811
rect 29 661 229 811
rect 287 661 487 811
rect -487 293 -287 443
rect -229 293 -29 443
rect 29 293 229 443
rect 287 293 487 443
rect -487 -75 -287 75
rect -229 -75 -29 75
rect 29 -75 229 75
rect 287 -75 487 75
rect -487 -443 -287 -293
rect -229 -443 -29 -293
rect 29 -443 229 -293
rect 287 -443 487 -293
rect -487 -811 -287 -661
rect -229 -811 -29 -661
rect 29 -811 229 -661
rect 287 -811 487 -661
<< mvndiff >>
rect -545 799 -487 811
rect -545 673 -533 799
rect -499 673 -487 799
rect -545 661 -487 673
rect -287 799 -229 811
rect -287 673 -275 799
rect -241 673 -229 799
rect -287 661 -229 673
rect -29 799 29 811
rect -29 673 -17 799
rect 17 673 29 799
rect -29 661 29 673
rect 229 799 287 811
rect 229 673 241 799
rect 275 673 287 799
rect 229 661 287 673
rect 487 799 545 811
rect 487 673 499 799
rect 533 673 545 799
rect 487 661 545 673
rect -545 431 -487 443
rect -545 305 -533 431
rect -499 305 -487 431
rect -545 293 -487 305
rect -287 431 -229 443
rect -287 305 -275 431
rect -241 305 -229 431
rect -287 293 -229 305
rect -29 431 29 443
rect -29 305 -17 431
rect 17 305 29 431
rect -29 293 29 305
rect 229 431 287 443
rect 229 305 241 431
rect 275 305 287 431
rect 229 293 287 305
rect 487 431 545 443
rect 487 305 499 431
rect 533 305 545 431
rect 487 293 545 305
rect -545 63 -487 75
rect -545 -63 -533 63
rect -499 -63 -487 63
rect -545 -75 -487 -63
rect -287 63 -229 75
rect -287 -63 -275 63
rect -241 -63 -229 63
rect -287 -75 -229 -63
rect -29 63 29 75
rect -29 -63 -17 63
rect 17 -63 29 63
rect -29 -75 29 -63
rect 229 63 287 75
rect 229 -63 241 63
rect 275 -63 287 63
rect 229 -75 287 -63
rect 487 63 545 75
rect 487 -63 499 63
rect 533 -63 545 63
rect 487 -75 545 -63
rect -545 -305 -487 -293
rect -545 -431 -533 -305
rect -499 -431 -487 -305
rect -545 -443 -487 -431
rect -287 -305 -229 -293
rect -287 -431 -275 -305
rect -241 -431 -229 -305
rect -287 -443 -229 -431
rect -29 -305 29 -293
rect -29 -431 -17 -305
rect 17 -431 29 -305
rect -29 -443 29 -431
rect 229 -305 287 -293
rect 229 -431 241 -305
rect 275 -431 287 -305
rect 229 -443 287 -431
rect 487 -305 545 -293
rect 487 -431 499 -305
rect 533 -431 545 -305
rect 487 -443 545 -431
rect -545 -673 -487 -661
rect -545 -799 -533 -673
rect -499 -799 -487 -673
rect -545 -811 -487 -799
rect -287 -673 -229 -661
rect -287 -799 -275 -673
rect -241 -799 -229 -673
rect -287 -811 -229 -799
rect -29 -673 29 -661
rect -29 -799 -17 -673
rect 17 -799 29 -673
rect -29 -811 29 -799
rect 229 -673 287 -661
rect 229 -799 241 -673
rect 275 -799 287 -673
rect 229 -811 287 -799
rect 487 -673 545 -661
rect 487 -799 499 -673
rect 533 -799 545 -673
rect 487 -811 545 -799
<< mvndiffc >>
rect -533 673 -499 799
rect -275 673 -241 799
rect -17 673 17 799
rect 241 673 275 799
rect 499 673 533 799
rect -533 305 -499 431
rect -275 305 -241 431
rect -17 305 17 431
rect 241 305 275 431
rect 499 305 533 431
rect -533 -63 -499 63
rect -275 -63 -241 63
rect -17 -63 17 63
rect 241 -63 275 63
rect 499 -63 533 63
rect -533 -431 -499 -305
rect -275 -431 -241 -305
rect -17 -431 17 -305
rect 241 -431 275 -305
rect 499 -431 533 -305
rect -533 -799 -499 -673
rect -275 -799 -241 -673
rect -17 -799 17 -673
rect 241 -799 275 -673
rect 499 -799 533 -673
<< mvpsubdiff >>
rect -679 1021 679 1033
rect -679 987 -571 1021
rect 571 987 679 1021
rect -679 975 679 987
rect -679 925 -621 975
rect -679 -925 -667 925
rect -633 -925 -621 925
rect 621 925 679 975
rect -679 -975 -621 -925
rect 621 -925 633 925
rect 667 -925 679 925
rect 621 -975 679 -925
rect -679 -987 679 -975
rect -679 -1021 -571 -987
rect 571 -1021 679 -987
rect -679 -1033 679 -1021
<< mvpsubdiffcont >>
rect -571 987 571 1021
rect -667 -925 -633 925
rect 633 -925 667 925
rect -571 -1021 571 -987
<< poly >>
rect -487 883 -287 899
rect -487 849 -471 883
rect -303 849 -287 883
rect -487 811 -287 849
rect -229 883 -29 899
rect -229 849 -213 883
rect -45 849 -29 883
rect -229 811 -29 849
rect 29 883 229 899
rect 29 849 45 883
rect 213 849 229 883
rect 29 811 229 849
rect 287 883 487 899
rect 287 849 303 883
rect 471 849 487 883
rect 287 811 487 849
rect -487 623 -287 661
rect -487 589 -471 623
rect -303 589 -287 623
rect -487 573 -287 589
rect -229 623 -29 661
rect -229 589 -213 623
rect -45 589 -29 623
rect -229 573 -29 589
rect 29 623 229 661
rect 29 589 45 623
rect 213 589 229 623
rect 29 573 229 589
rect 287 623 487 661
rect 287 589 303 623
rect 471 589 487 623
rect 287 573 487 589
rect -487 515 -287 531
rect -487 481 -471 515
rect -303 481 -287 515
rect -487 443 -287 481
rect -229 515 -29 531
rect -229 481 -213 515
rect -45 481 -29 515
rect -229 443 -29 481
rect 29 515 229 531
rect 29 481 45 515
rect 213 481 229 515
rect 29 443 229 481
rect 287 515 487 531
rect 287 481 303 515
rect 471 481 487 515
rect 287 443 487 481
rect -487 255 -287 293
rect -487 221 -471 255
rect -303 221 -287 255
rect -487 205 -287 221
rect -229 255 -29 293
rect -229 221 -213 255
rect -45 221 -29 255
rect -229 205 -29 221
rect 29 255 229 293
rect 29 221 45 255
rect 213 221 229 255
rect 29 205 229 221
rect 287 255 487 293
rect 287 221 303 255
rect 471 221 487 255
rect 287 205 487 221
rect -487 147 -287 163
rect -487 113 -471 147
rect -303 113 -287 147
rect -487 75 -287 113
rect -229 147 -29 163
rect -229 113 -213 147
rect -45 113 -29 147
rect -229 75 -29 113
rect 29 147 229 163
rect 29 113 45 147
rect 213 113 229 147
rect 29 75 229 113
rect 287 147 487 163
rect 287 113 303 147
rect 471 113 487 147
rect 287 75 487 113
rect -487 -113 -287 -75
rect -487 -147 -471 -113
rect -303 -147 -287 -113
rect -487 -163 -287 -147
rect -229 -113 -29 -75
rect -229 -147 -213 -113
rect -45 -147 -29 -113
rect -229 -163 -29 -147
rect 29 -113 229 -75
rect 29 -147 45 -113
rect 213 -147 229 -113
rect 29 -163 229 -147
rect 287 -113 487 -75
rect 287 -147 303 -113
rect 471 -147 487 -113
rect 287 -163 487 -147
rect -487 -221 -287 -205
rect -487 -255 -471 -221
rect -303 -255 -287 -221
rect -487 -293 -287 -255
rect -229 -221 -29 -205
rect -229 -255 -213 -221
rect -45 -255 -29 -221
rect -229 -293 -29 -255
rect 29 -221 229 -205
rect 29 -255 45 -221
rect 213 -255 229 -221
rect 29 -293 229 -255
rect 287 -221 487 -205
rect 287 -255 303 -221
rect 471 -255 487 -221
rect 287 -293 487 -255
rect -487 -481 -287 -443
rect -487 -515 -471 -481
rect -303 -515 -287 -481
rect -487 -531 -287 -515
rect -229 -481 -29 -443
rect -229 -515 -213 -481
rect -45 -515 -29 -481
rect -229 -531 -29 -515
rect 29 -481 229 -443
rect 29 -515 45 -481
rect 213 -515 229 -481
rect 29 -531 229 -515
rect 287 -481 487 -443
rect 287 -515 303 -481
rect 471 -515 487 -481
rect 287 -531 487 -515
rect -487 -589 -287 -573
rect -487 -623 -471 -589
rect -303 -623 -287 -589
rect -487 -661 -287 -623
rect -229 -589 -29 -573
rect -229 -623 -213 -589
rect -45 -623 -29 -589
rect -229 -661 -29 -623
rect 29 -589 229 -573
rect 29 -623 45 -589
rect 213 -623 229 -589
rect 29 -661 229 -623
rect 287 -589 487 -573
rect 287 -623 303 -589
rect 471 -623 487 -589
rect 287 -661 487 -623
rect -487 -849 -287 -811
rect -487 -883 -471 -849
rect -303 -883 -287 -849
rect -487 -899 -287 -883
rect -229 -849 -29 -811
rect -229 -883 -213 -849
rect -45 -883 -29 -849
rect -229 -899 -29 -883
rect 29 -849 229 -811
rect 29 -883 45 -849
rect 213 -883 229 -849
rect 29 -899 229 -883
rect 287 -849 487 -811
rect 287 -883 303 -849
rect 471 -883 487 -849
rect 287 -899 487 -883
<< polycont >>
rect -471 849 -303 883
rect -213 849 -45 883
rect 45 849 213 883
rect 303 849 471 883
rect -471 589 -303 623
rect -213 589 -45 623
rect 45 589 213 623
rect 303 589 471 623
rect -471 481 -303 515
rect -213 481 -45 515
rect 45 481 213 515
rect 303 481 471 515
rect -471 221 -303 255
rect -213 221 -45 255
rect 45 221 213 255
rect 303 221 471 255
rect -471 113 -303 147
rect -213 113 -45 147
rect 45 113 213 147
rect 303 113 471 147
rect -471 -147 -303 -113
rect -213 -147 -45 -113
rect 45 -147 213 -113
rect 303 -147 471 -113
rect -471 -255 -303 -221
rect -213 -255 -45 -221
rect 45 -255 213 -221
rect 303 -255 471 -221
rect -471 -515 -303 -481
rect -213 -515 -45 -481
rect 45 -515 213 -481
rect 303 -515 471 -481
rect -471 -623 -303 -589
rect -213 -623 -45 -589
rect 45 -623 213 -589
rect 303 -623 471 -589
rect -471 -883 -303 -849
rect -213 -883 -45 -849
rect 45 -883 213 -849
rect 303 -883 471 -849
<< locali >>
rect -667 987 -571 1021
rect 571 987 667 1021
rect -667 925 -633 987
rect 633 925 667 987
rect -487 849 -471 883
rect -303 849 -287 883
rect -229 849 -213 883
rect -45 849 -29 883
rect 29 849 45 883
rect 213 849 229 883
rect 287 849 303 883
rect 471 849 487 883
rect -533 799 -499 815
rect -533 657 -499 673
rect -275 799 -241 815
rect -275 657 -241 673
rect -17 799 17 815
rect -17 657 17 673
rect 241 799 275 815
rect 241 657 275 673
rect 499 799 533 815
rect 499 657 533 673
rect -487 589 -471 623
rect -303 589 -287 623
rect -229 589 -213 623
rect -45 589 -29 623
rect 29 589 45 623
rect 213 589 229 623
rect 287 589 303 623
rect 471 589 487 623
rect -487 481 -471 515
rect -303 481 -287 515
rect -229 481 -213 515
rect -45 481 -29 515
rect 29 481 45 515
rect 213 481 229 515
rect 287 481 303 515
rect 471 481 487 515
rect -533 431 -499 447
rect -533 289 -499 305
rect -275 431 -241 447
rect -275 289 -241 305
rect -17 431 17 447
rect -17 289 17 305
rect 241 431 275 447
rect 241 289 275 305
rect 499 431 533 447
rect 499 289 533 305
rect -487 221 -471 255
rect -303 221 -287 255
rect -229 221 -213 255
rect -45 221 -29 255
rect 29 221 45 255
rect 213 221 229 255
rect 287 221 303 255
rect 471 221 487 255
rect -487 113 -471 147
rect -303 113 -287 147
rect -229 113 -213 147
rect -45 113 -29 147
rect 29 113 45 147
rect 213 113 229 147
rect 287 113 303 147
rect 471 113 487 147
rect -533 63 -499 79
rect -533 -79 -499 -63
rect -275 63 -241 79
rect -275 -79 -241 -63
rect -17 63 17 79
rect -17 -79 17 -63
rect 241 63 275 79
rect 241 -79 275 -63
rect 499 63 533 79
rect 499 -79 533 -63
rect -487 -147 -471 -113
rect -303 -147 -287 -113
rect -229 -147 -213 -113
rect -45 -147 -29 -113
rect 29 -147 45 -113
rect 213 -147 229 -113
rect 287 -147 303 -113
rect 471 -147 487 -113
rect -487 -255 -471 -221
rect -303 -255 -287 -221
rect -229 -255 -213 -221
rect -45 -255 -29 -221
rect 29 -255 45 -221
rect 213 -255 229 -221
rect 287 -255 303 -221
rect 471 -255 487 -221
rect -533 -305 -499 -289
rect -533 -447 -499 -431
rect -275 -305 -241 -289
rect -275 -447 -241 -431
rect -17 -305 17 -289
rect -17 -447 17 -431
rect 241 -305 275 -289
rect 241 -447 275 -431
rect 499 -305 533 -289
rect 499 -447 533 -431
rect -487 -515 -471 -481
rect -303 -515 -287 -481
rect -229 -515 -213 -481
rect -45 -515 -29 -481
rect 29 -515 45 -481
rect 213 -515 229 -481
rect 287 -515 303 -481
rect 471 -515 487 -481
rect -487 -623 -471 -589
rect -303 -623 -287 -589
rect -229 -623 -213 -589
rect -45 -623 -29 -589
rect 29 -623 45 -589
rect 213 -623 229 -589
rect 287 -623 303 -589
rect 471 -623 487 -589
rect -533 -673 -499 -657
rect -533 -815 -499 -799
rect -275 -673 -241 -657
rect -275 -815 -241 -799
rect -17 -673 17 -657
rect -17 -815 17 -799
rect 241 -673 275 -657
rect 241 -815 275 -799
rect 499 -673 533 -657
rect 499 -815 533 -799
rect -487 -883 -471 -849
rect -303 -883 -287 -849
rect -229 -883 -213 -849
rect -45 -883 -29 -849
rect 29 -883 45 -849
rect 213 -883 229 -849
rect 287 -883 303 -849
rect 471 -883 487 -849
rect -667 -987 -633 -925
rect 633 -987 667 -925
rect -667 -1021 -571 -987
rect 571 -1021 667 -987
<< viali >>
rect -471 849 -303 883
rect -213 849 -45 883
rect 45 849 213 883
rect 303 849 471 883
rect -533 673 -499 799
rect -275 673 -241 799
rect -17 673 17 799
rect 241 673 275 799
rect 499 673 533 799
rect -471 589 -303 623
rect -213 589 -45 623
rect 45 589 213 623
rect 303 589 471 623
rect -471 481 -303 515
rect -213 481 -45 515
rect 45 481 213 515
rect 303 481 471 515
rect -533 305 -499 431
rect -275 305 -241 431
rect -17 305 17 431
rect 241 305 275 431
rect 499 305 533 431
rect -471 221 -303 255
rect -213 221 -45 255
rect 45 221 213 255
rect 303 221 471 255
rect -471 113 -303 147
rect -213 113 -45 147
rect 45 113 213 147
rect 303 113 471 147
rect -533 -63 -499 63
rect -275 -63 -241 63
rect -17 -63 17 63
rect 241 -63 275 63
rect 499 -63 533 63
rect -471 -147 -303 -113
rect -213 -147 -45 -113
rect 45 -147 213 -113
rect 303 -147 471 -113
rect -471 -255 -303 -221
rect -213 -255 -45 -221
rect 45 -255 213 -221
rect 303 -255 471 -221
rect -533 -431 -499 -305
rect -275 -431 -241 -305
rect -17 -431 17 -305
rect 241 -431 275 -305
rect 499 -431 533 -305
rect -471 -515 -303 -481
rect -213 -515 -45 -481
rect 45 -515 213 -481
rect 303 -515 471 -481
rect -471 -623 -303 -589
rect -213 -623 -45 -589
rect 45 -623 213 -589
rect 303 -623 471 -589
rect -533 -799 -499 -673
rect -275 -799 -241 -673
rect -17 -799 17 -673
rect 241 -799 275 -673
rect 499 -799 533 -673
rect -471 -883 -303 -849
rect -213 -883 -45 -849
rect 45 -883 213 -849
rect 303 -883 471 -849
<< metal1 >>
rect -483 883 -291 889
rect -483 849 -471 883
rect -303 849 -291 883
rect -483 843 -291 849
rect -225 883 -33 889
rect -225 849 -213 883
rect -45 849 -33 883
rect -225 843 -33 849
rect 33 883 225 889
rect 33 849 45 883
rect 213 849 225 883
rect 33 843 225 849
rect 291 883 483 889
rect 291 849 303 883
rect 471 849 483 883
rect 291 843 483 849
rect -539 799 -493 811
rect -539 673 -533 799
rect -499 673 -493 799
rect -539 661 -493 673
rect -281 799 -235 811
rect -281 673 -275 799
rect -241 673 -235 799
rect -281 661 -235 673
rect -23 799 23 811
rect -23 673 -17 799
rect 17 673 23 799
rect -23 661 23 673
rect 235 799 281 811
rect 235 673 241 799
rect 275 673 281 799
rect 235 661 281 673
rect 493 799 539 811
rect 493 673 499 799
rect 533 673 539 799
rect 493 661 539 673
rect -483 623 -291 629
rect -483 589 -471 623
rect -303 589 -291 623
rect -483 583 -291 589
rect -225 623 -33 629
rect -225 589 -213 623
rect -45 589 -33 623
rect -225 583 -33 589
rect 33 623 225 629
rect 33 589 45 623
rect 213 589 225 623
rect 33 583 225 589
rect 291 623 483 629
rect 291 589 303 623
rect 471 589 483 623
rect 291 583 483 589
rect -483 515 -291 521
rect -483 481 -471 515
rect -303 481 -291 515
rect -483 475 -291 481
rect -225 515 -33 521
rect -225 481 -213 515
rect -45 481 -33 515
rect -225 475 -33 481
rect 33 515 225 521
rect 33 481 45 515
rect 213 481 225 515
rect 33 475 225 481
rect 291 515 483 521
rect 291 481 303 515
rect 471 481 483 515
rect 291 475 483 481
rect -539 431 -493 443
rect -539 305 -533 431
rect -499 305 -493 431
rect -539 293 -493 305
rect -281 431 -235 443
rect -281 305 -275 431
rect -241 305 -235 431
rect -281 293 -235 305
rect -23 431 23 443
rect -23 305 -17 431
rect 17 305 23 431
rect -23 293 23 305
rect 235 431 281 443
rect 235 305 241 431
rect 275 305 281 431
rect 235 293 281 305
rect 493 431 539 443
rect 493 305 499 431
rect 533 305 539 431
rect 493 293 539 305
rect -483 255 -291 261
rect -483 221 -471 255
rect -303 221 -291 255
rect -483 215 -291 221
rect -225 255 -33 261
rect -225 221 -213 255
rect -45 221 -33 255
rect -225 215 -33 221
rect 33 255 225 261
rect 33 221 45 255
rect 213 221 225 255
rect 33 215 225 221
rect 291 255 483 261
rect 291 221 303 255
rect 471 221 483 255
rect 291 215 483 221
rect -483 147 -291 153
rect -483 113 -471 147
rect -303 113 -291 147
rect -483 107 -291 113
rect -225 147 -33 153
rect -225 113 -213 147
rect -45 113 -33 147
rect -225 107 -33 113
rect 33 147 225 153
rect 33 113 45 147
rect 213 113 225 147
rect 33 107 225 113
rect 291 147 483 153
rect 291 113 303 147
rect 471 113 483 147
rect 291 107 483 113
rect -539 63 -493 75
rect -539 -63 -533 63
rect -499 -63 -493 63
rect -539 -75 -493 -63
rect -281 63 -235 75
rect -281 -63 -275 63
rect -241 -63 -235 63
rect -281 -75 -235 -63
rect -23 63 23 75
rect -23 -63 -17 63
rect 17 -63 23 63
rect -23 -75 23 -63
rect 235 63 281 75
rect 235 -63 241 63
rect 275 -63 281 63
rect 235 -75 281 -63
rect 493 63 539 75
rect 493 -63 499 63
rect 533 -63 539 63
rect 493 -75 539 -63
rect -483 -113 -291 -107
rect -483 -147 -471 -113
rect -303 -147 -291 -113
rect -483 -153 -291 -147
rect -225 -113 -33 -107
rect -225 -147 -213 -113
rect -45 -147 -33 -113
rect -225 -153 -33 -147
rect 33 -113 225 -107
rect 33 -147 45 -113
rect 213 -147 225 -113
rect 33 -153 225 -147
rect 291 -113 483 -107
rect 291 -147 303 -113
rect 471 -147 483 -113
rect 291 -153 483 -147
rect -483 -221 -291 -215
rect -483 -255 -471 -221
rect -303 -255 -291 -221
rect -483 -261 -291 -255
rect -225 -221 -33 -215
rect -225 -255 -213 -221
rect -45 -255 -33 -221
rect -225 -261 -33 -255
rect 33 -221 225 -215
rect 33 -255 45 -221
rect 213 -255 225 -221
rect 33 -261 225 -255
rect 291 -221 483 -215
rect 291 -255 303 -221
rect 471 -255 483 -221
rect 291 -261 483 -255
rect -539 -305 -493 -293
rect -539 -431 -533 -305
rect -499 -431 -493 -305
rect -539 -443 -493 -431
rect -281 -305 -235 -293
rect -281 -431 -275 -305
rect -241 -431 -235 -305
rect -281 -443 -235 -431
rect -23 -305 23 -293
rect -23 -431 -17 -305
rect 17 -431 23 -305
rect -23 -443 23 -431
rect 235 -305 281 -293
rect 235 -431 241 -305
rect 275 -431 281 -305
rect 235 -443 281 -431
rect 493 -305 539 -293
rect 493 -431 499 -305
rect 533 -431 539 -305
rect 493 -443 539 -431
rect -483 -481 -291 -475
rect -483 -515 -471 -481
rect -303 -515 -291 -481
rect -483 -521 -291 -515
rect -225 -481 -33 -475
rect -225 -515 -213 -481
rect -45 -515 -33 -481
rect -225 -521 -33 -515
rect 33 -481 225 -475
rect 33 -515 45 -481
rect 213 -515 225 -481
rect 33 -521 225 -515
rect 291 -481 483 -475
rect 291 -515 303 -481
rect 471 -515 483 -481
rect 291 -521 483 -515
rect -483 -589 -291 -583
rect -483 -623 -471 -589
rect -303 -623 -291 -589
rect -483 -629 -291 -623
rect -225 -589 -33 -583
rect -225 -623 -213 -589
rect -45 -623 -33 -589
rect -225 -629 -33 -623
rect 33 -589 225 -583
rect 33 -623 45 -589
rect 213 -623 225 -589
rect 33 -629 225 -623
rect 291 -589 483 -583
rect 291 -623 303 -589
rect 471 -623 483 -589
rect 291 -629 483 -623
rect -539 -673 -493 -661
rect -539 -799 -533 -673
rect -499 -799 -493 -673
rect -539 -811 -493 -799
rect -281 -673 -235 -661
rect -281 -799 -275 -673
rect -241 -799 -235 -673
rect -281 -811 -235 -799
rect -23 -673 23 -661
rect -23 -799 -17 -673
rect 17 -799 23 -673
rect -23 -811 23 -799
rect 235 -673 281 -661
rect 235 -799 241 -673
rect 275 -799 281 -673
rect 235 -811 281 -799
rect 493 -673 539 -661
rect 493 -799 499 -673
rect 533 -799 539 -673
rect 493 -811 539 -799
rect -483 -849 -291 -843
rect -483 -883 -471 -849
rect -303 -883 -291 -849
rect -483 -889 -291 -883
rect -225 -849 -33 -843
rect -225 -883 -213 -849
rect -45 -883 -33 -849
rect -225 -889 -33 -883
rect 33 -849 225 -843
rect 33 -883 45 -849
rect 213 -883 225 -849
rect 33 -889 225 -883
rect 291 -849 483 -843
rect 291 -883 303 -849
rect 471 -883 483 -849
rect 291 -889 483 -883
<< properties >>
string FIXED_BBOX -650 -1004 650 1004
string gencell sky130_fd_pr__nfet_g5v0d10v5
string library sky130
string parameters w 0.75 l 1.0 m 5 nf 4 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
