magic
tech sky130A
magscale 1 2
timestamp 1716807968
<< pwell >>
rect -328 -10329 328 10329
<< mvnmos >>
rect -100 9271 100 10071
rect -100 8253 100 9053
rect -100 7235 100 8035
rect -100 6217 100 7017
rect -100 5199 100 5999
rect -100 4181 100 4981
rect -100 3163 100 3963
rect -100 2145 100 2945
rect -100 1127 100 1927
rect -100 109 100 909
rect -100 -909 100 -109
rect -100 -1927 100 -1127
rect -100 -2945 100 -2145
rect -100 -3963 100 -3163
rect -100 -4981 100 -4181
rect -100 -5999 100 -5199
rect -100 -7017 100 -6217
rect -100 -8035 100 -7235
rect -100 -9053 100 -8253
rect -100 -10071 100 -9271
<< mvndiff >>
rect -158 10059 -100 10071
rect -158 9283 -146 10059
rect -112 9283 -100 10059
rect -158 9271 -100 9283
rect 100 10059 158 10071
rect 100 9283 112 10059
rect 146 9283 158 10059
rect 100 9271 158 9283
rect -158 9041 -100 9053
rect -158 8265 -146 9041
rect -112 8265 -100 9041
rect -158 8253 -100 8265
rect 100 9041 158 9053
rect 100 8265 112 9041
rect 146 8265 158 9041
rect 100 8253 158 8265
rect -158 8023 -100 8035
rect -158 7247 -146 8023
rect -112 7247 -100 8023
rect -158 7235 -100 7247
rect 100 8023 158 8035
rect 100 7247 112 8023
rect 146 7247 158 8023
rect 100 7235 158 7247
rect -158 7005 -100 7017
rect -158 6229 -146 7005
rect -112 6229 -100 7005
rect -158 6217 -100 6229
rect 100 7005 158 7017
rect 100 6229 112 7005
rect 146 6229 158 7005
rect 100 6217 158 6229
rect -158 5987 -100 5999
rect -158 5211 -146 5987
rect -112 5211 -100 5987
rect -158 5199 -100 5211
rect 100 5987 158 5999
rect 100 5211 112 5987
rect 146 5211 158 5987
rect 100 5199 158 5211
rect -158 4969 -100 4981
rect -158 4193 -146 4969
rect -112 4193 -100 4969
rect -158 4181 -100 4193
rect 100 4969 158 4981
rect 100 4193 112 4969
rect 146 4193 158 4969
rect 100 4181 158 4193
rect -158 3951 -100 3963
rect -158 3175 -146 3951
rect -112 3175 -100 3951
rect -158 3163 -100 3175
rect 100 3951 158 3963
rect 100 3175 112 3951
rect 146 3175 158 3951
rect 100 3163 158 3175
rect -158 2933 -100 2945
rect -158 2157 -146 2933
rect -112 2157 -100 2933
rect -158 2145 -100 2157
rect 100 2933 158 2945
rect 100 2157 112 2933
rect 146 2157 158 2933
rect 100 2145 158 2157
rect -158 1915 -100 1927
rect -158 1139 -146 1915
rect -112 1139 -100 1915
rect -158 1127 -100 1139
rect 100 1915 158 1927
rect 100 1139 112 1915
rect 146 1139 158 1915
rect 100 1127 158 1139
rect -158 897 -100 909
rect -158 121 -146 897
rect -112 121 -100 897
rect -158 109 -100 121
rect 100 897 158 909
rect 100 121 112 897
rect 146 121 158 897
rect 100 109 158 121
rect -158 -121 -100 -109
rect -158 -897 -146 -121
rect -112 -897 -100 -121
rect -158 -909 -100 -897
rect 100 -121 158 -109
rect 100 -897 112 -121
rect 146 -897 158 -121
rect 100 -909 158 -897
rect -158 -1139 -100 -1127
rect -158 -1915 -146 -1139
rect -112 -1915 -100 -1139
rect -158 -1927 -100 -1915
rect 100 -1139 158 -1127
rect 100 -1915 112 -1139
rect 146 -1915 158 -1139
rect 100 -1927 158 -1915
rect -158 -2157 -100 -2145
rect -158 -2933 -146 -2157
rect -112 -2933 -100 -2157
rect -158 -2945 -100 -2933
rect 100 -2157 158 -2145
rect 100 -2933 112 -2157
rect 146 -2933 158 -2157
rect 100 -2945 158 -2933
rect -158 -3175 -100 -3163
rect -158 -3951 -146 -3175
rect -112 -3951 -100 -3175
rect -158 -3963 -100 -3951
rect 100 -3175 158 -3163
rect 100 -3951 112 -3175
rect 146 -3951 158 -3175
rect 100 -3963 158 -3951
rect -158 -4193 -100 -4181
rect -158 -4969 -146 -4193
rect -112 -4969 -100 -4193
rect -158 -4981 -100 -4969
rect 100 -4193 158 -4181
rect 100 -4969 112 -4193
rect 146 -4969 158 -4193
rect 100 -4981 158 -4969
rect -158 -5211 -100 -5199
rect -158 -5987 -146 -5211
rect -112 -5987 -100 -5211
rect -158 -5999 -100 -5987
rect 100 -5211 158 -5199
rect 100 -5987 112 -5211
rect 146 -5987 158 -5211
rect 100 -5999 158 -5987
rect -158 -6229 -100 -6217
rect -158 -7005 -146 -6229
rect -112 -7005 -100 -6229
rect -158 -7017 -100 -7005
rect 100 -6229 158 -6217
rect 100 -7005 112 -6229
rect 146 -7005 158 -6229
rect 100 -7017 158 -7005
rect -158 -7247 -100 -7235
rect -158 -8023 -146 -7247
rect -112 -8023 -100 -7247
rect -158 -8035 -100 -8023
rect 100 -7247 158 -7235
rect 100 -8023 112 -7247
rect 146 -8023 158 -7247
rect 100 -8035 158 -8023
rect -158 -8265 -100 -8253
rect -158 -9041 -146 -8265
rect -112 -9041 -100 -8265
rect -158 -9053 -100 -9041
rect 100 -8265 158 -8253
rect 100 -9041 112 -8265
rect 146 -9041 158 -8265
rect 100 -9053 158 -9041
rect -158 -9283 -100 -9271
rect -158 -10059 -146 -9283
rect -112 -10059 -100 -9283
rect -158 -10071 -100 -10059
rect 100 -9283 158 -9271
rect 100 -10059 112 -9283
rect 146 -10059 158 -9283
rect 100 -10071 158 -10059
<< mvndiffc >>
rect -146 9283 -112 10059
rect 112 9283 146 10059
rect -146 8265 -112 9041
rect 112 8265 146 9041
rect -146 7247 -112 8023
rect 112 7247 146 8023
rect -146 6229 -112 7005
rect 112 6229 146 7005
rect -146 5211 -112 5987
rect 112 5211 146 5987
rect -146 4193 -112 4969
rect 112 4193 146 4969
rect -146 3175 -112 3951
rect 112 3175 146 3951
rect -146 2157 -112 2933
rect 112 2157 146 2933
rect -146 1139 -112 1915
rect 112 1139 146 1915
rect -146 121 -112 897
rect 112 121 146 897
rect -146 -897 -112 -121
rect 112 -897 146 -121
rect -146 -1915 -112 -1139
rect 112 -1915 146 -1139
rect -146 -2933 -112 -2157
rect 112 -2933 146 -2157
rect -146 -3951 -112 -3175
rect 112 -3951 146 -3175
rect -146 -4969 -112 -4193
rect 112 -4969 146 -4193
rect -146 -5987 -112 -5211
rect 112 -5987 146 -5211
rect -146 -7005 -112 -6229
rect 112 -7005 146 -6229
rect -146 -8023 -112 -7247
rect 112 -8023 146 -7247
rect -146 -9041 -112 -8265
rect 112 -9041 146 -8265
rect -146 -10059 -112 -9283
rect 112 -10059 146 -9283
<< mvpsubdiff >>
rect -292 10281 292 10293
rect -292 10247 -184 10281
rect 184 10247 292 10281
rect -292 10235 292 10247
rect -292 10185 -234 10235
rect -292 -10185 -280 10185
rect -246 -10185 -234 10185
rect 234 10185 292 10235
rect -292 -10235 -234 -10185
rect 234 -10185 246 10185
rect 280 -10185 292 10185
rect 234 -10235 292 -10185
rect -292 -10247 292 -10235
rect -292 -10281 -184 -10247
rect 184 -10281 292 -10247
rect -292 -10293 292 -10281
<< mvpsubdiffcont >>
rect -184 10247 184 10281
rect -280 -10185 -246 10185
rect 246 -10185 280 10185
rect -184 -10281 184 -10247
<< poly >>
rect -100 10143 100 10159
rect -100 10109 -84 10143
rect 84 10109 100 10143
rect -100 10071 100 10109
rect -100 9233 100 9271
rect -100 9199 -84 9233
rect 84 9199 100 9233
rect -100 9183 100 9199
rect -100 9125 100 9141
rect -100 9091 -84 9125
rect 84 9091 100 9125
rect -100 9053 100 9091
rect -100 8215 100 8253
rect -100 8181 -84 8215
rect 84 8181 100 8215
rect -100 8165 100 8181
rect -100 8107 100 8123
rect -100 8073 -84 8107
rect 84 8073 100 8107
rect -100 8035 100 8073
rect -100 7197 100 7235
rect -100 7163 -84 7197
rect 84 7163 100 7197
rect -100 7147 100 7163
rect -100 7089 100 7105
rect -100 7055 -84 7089
rect 84 7055 100 7089
rect -100 7017 100 7055
rect -100 6179 100 6217
rect -100 6145 -84 6179
rect 84 6145 100 6179
rect -100 6129 100 6145
rect -100 6071 100 6087
rect -100 6037 -84 6071
rect 84 6037 100 6071
rect -100 5999 100 6037
rect -100 5161 100 5199
rect -100 5127 -84 5161
rect 84 5127 100 5161
rect -100 5111 100 5127
rect -100 5053 100 5069
rect -100 5019 -84 5053
rect 84 5019 100 5053
rect -100 4981 100 5019
rect -100 4143 100 4181
rect -100 4109 -84 4143
rect 84 4109 100 4143
rect -100 4093 100 4109
rect -100 4035 100 4051
rect -100 4001 -84 4035
rect 84 4001 100 4035
rect -100 3963 100 4001
rect -100 3125 100 3163
rect -100 3091 -84 3125
rect 84 3091 100 3125
rect -100 3075 100 3091
rect -100 3017 100 3033
rect -100 2983 -84 3017
rect 84 2983 100 3017
rect -100 2945 100 2983
rect -100 2107 100 2145
rect -100 2073 -84 2107
rect 84 2073 100 2107
rect -100 2057 100 2073
rect -100 1999 100 2015
rect -100 1965 -84 1999
rect 84 1965 100 1999
rect -100 1927 100 1965
rect -100 1089 100 1127
rect -100 1055 -84 1089
rect 84 1055 100 1089
rect -100 1039 100 1055
rect -100 981 100 997
rect -100 947 -84 981
rect 84 947 100 981
rect -100 909 100 947
rect -100 71 100 109
rect -100 37 -84 71
rect 84 37 100 71
rect -100 21 100 37
rect -100 -37 100 -21
rect -100 -71 -84 -37
rect 84 -71 100 -37
rect -100 -109 100 -71
rect -100 -947 100 -909
rect -100 -981 -84 -947
rect 84 -981 100 -947
rect -100 -997 100 -981
rect -100 -1055 100 -1039
rect -100 -1089 -84 -1055
rect 84 -1089 100 -1055
rect -100 -1127 100 -1089
rect -100 -1965 100 -1927
rect -100 -1999 -84 -1965
rect 84 -1999 100 -1965
rect -100 -2015 100 -1999
rect -100 -2073 100 -2057
rect -100 -2107 -84 -2073
rect 84 -2107 100 -2073
rect -100 -2145 100 -2107
rect -100 -2983 100 -2945
rect -100 -3017 -84 -2983
rect 84 -3017 100 -2983
rect -100 -3033 100 -3017
rect -100 -3091 100 -3075
rect -100 -3125 -84 -3091
rect 84 -3125 100 -3091
rect -100 -3163 100 -3125
rect -100 -4001 100 -3963
rect -100 -4035 -84 -4001
rect 84 -4035 100 -4001
rect -100 -4051 100 -4035
rect -100 -4109 100 -4093
rect -100 -4143 -84 -4109
rect 84 -4143 100 -4109
rect -100 -4181 100 -4143
rect -100 -5019 100 -4981
rect -100 -5053 -84 -5019
rect 84 -5053 100 -5019
rect -100 -5069 100 -5053
rect -100 -5127 100 -5111
rect -100 -5161 -84 -5127
rect 84 -5161 100 -5127
rect -100 -5199 100 -5161
rect -100 -6037 100 -5999
rect -100 -6071 -84 -6037
rect 84 -6071 100 -6037
rect -100 -6087 100 -6071
rect -100 -6145 100 -6129
rect -100 -6179 -84 -6145
rect 84 -6179 100 -6145
rect -100 -6217 100 -6179
rect -100 -7055 100 -7017
rect -100 -7089 -84 -7055
rect 84 -7089 100 -7055
rect -100 -7105 100 -7089
rect -100 -7163 100 -7147
rect -100 -7197 -84 -7163
rect 84 -7197 100 -7163
rect -100 -7235 100 -7197
rect -100 -8073 100 -8035
rect -100 -8107 -84 -8073
rect 84 -8107 100 -8073
rect -100 -8123 100 -8107
rect -100 -8181 100 -8165
rect -100 -8215 -84 -8181
rect 84 -8215 100 -8181
rect -100 -8253 100 -8215
rect -100 -9091 100 -9053
rect -100 -9125 -84 -9091
rect 84 -9125 100 -9091
rect -100 -9141 100 -9125
rect -100 -9199 100 -9183
rect -100 -9233 -84 -9199
rect 84 -9233 100 -9199
rect -100 -9271 100 -9233
rect -100 -10109 100 -10071
rect -100 -10143 -84 -10109
rect 84 -10143 100 -10109
rect -100 -10159 100 -10143
<< polycont >>
rect -84 10109 84 10143
rect -84 9199 84 9233
rect -84 9091 84 9125
rect -84 8181 84 8215
rect -84 8073 84 8107
rect -84 7163 84 7197
rect -84 7055 84 7089
rect -84 6145 84 6179
rect -84 6037 84 6071
rect -84 5127 84 5161
rect -84 5019 84 5053
rect -84 4109 84 4143
rect -84 4001 84 4035
rect -84 3091 84 3125
rect -84 2983 84 3017
rect -84 2073 84 2107
rect -84 1965 84 1999
rect -84 1055 84 1089
rect -84 947 84 981
rect -84 37 84 71
rect -84 -71 84 -37
rect -84 -981 84 -947
rect -84 -1089 84 -1055
rect -84 -1999 84 -1965
rect -84 -2107 84 -2073
rect -84 -3017 84 -2983
rect -84 -3125 84 -3091
rect -84 -4035 84 -4001
rect -84 -4143 84 -4109
rect -84 -5053 84 -5019
rect -84 -5161 84 -5127
rect -84 -6071 84 -6037
rect -84 -6179 84 -6145
rect -84 -7089 84 -7055
rect -84 -7197 84 -7163
rect -84 -8107 84 -8073
rect -84 -8215 84 -8181
rect -84 -9125 84 -9091
rect -84 -9233 84 -9199
rect -84 -10143 84 -10109
<< locali >>
rect -280 10247 -184 10281
rect 184 10247 280 10281
rect -280 10185 -246 10247
rect 246 10185 280 10247
rect -100 10109 -84 10143
rect 84 10109 100 10143
rect -146 10059 -112 10075
rect -146 9267 -112 9283
rect 112 10059 146 10075
rect 112 9267 146 9283
rect -100 9199 -84 9233
rect 84 9199 100 9233
rect -100 9091 -84 9125
rect 84 9091 100 9125
rect -146 9041 -112 9057
rect -146 8249 -112 8265
rect 112 9041 146 9057
rect 112 8249 146 8265
rect -100 8181 -84 8215
rect 84 8181 100 8215
rect -100 8073 -84 8107
rect 84 8073 100 8107
rect -146 8023 -112 8039
rect -146 7231 -112 7247
rect 112 8023 146 8039
rect 112 7231 146 7247
rect -100 7163 -84 7197
rect 84 7163 100 7197
rect -100 7055 -84 7089
rect 84 7055 100 7089
rect -146 7005 -112 7021
rect -146 6213 -112 6229
rect 112 7005 146 7021
rect 112 6213 146 6229
rect -100 6145 -84 6179
rect 84 6145 100 6179
rect -100 6037 -84 6071
rect 84 6037 100 6071
rect -146 5987 -112 6003
rect -146 5195 -112 5211
rect 112 5987 146 6003
rect 112 5195 146 5211
rect -100 5127 -84 5161
rect 84 5127 100 5161
rect -100 5019 -84 5053
rect 84 5019 100 5053
rect -146 4969 -112 4985
rect -146 4177 -112 4193
rect 112 4969 146 4985
rect 112 4177 146 4193
rect -100 4109 -84 4143
rect 84 4109 100 4143
rect -100 4001 -84 4035
rect 84 4001 100 4035
rect -146 3951 -112 3967
rect -146 3159 -112 3175
rect 112 3951 146 3967
rect 112 3159 146 3175
rect -100 3091 -84 3125
rect 84 3091 100 3125
rect -100 2983 -84 3017
rect 84 2983 100 3017
rect -146 2933 -112 2949
rect -146 2141 -112 2157
rect 112 2933 146 2949
rect 112 2141 146 2157
rect -100 2073 -84 2107
rect 84 2073 100 2107
rect -100 1965 -84 1999
rect 84 1965 100 1999
rect -146 1915 -112 1931
rect -146 1123 -112 1139
rect 112 1915 146 1931
rect 112 1123 146 1139
rect -100 1055 -84 1089
rect 84 1055 100 1089
rect -100 947 -84 981
rect 84 947 100 981
rect -146 897 -112 913
rect -146 105 -112 121
rect 112 897 146 913
rect 112 105 146 121
rect -100 37 -84 71
rect 84 37 100 71
rect -100 -71 -84 -37
rect 84 -71 100 -37
rect -146 -121 -112 -105
rect -146 -913 -112 -897
rect 112 -121 146 -105
rect 112 -913 146 -897
rect -100 -981 -84 -947
rect 84 -981 100 -947
rect -100 -1089 -84 -1055
rect 84 -1089 100 -1055
rect -146 -1139 -112 -1123
rect -146 -1931 -112 -1915
rect 112 -1139 146 -1123
rect 112 -1931 146 -1915
rect -100 -1999 -84 -1965
rect 84 -1999 100 -1965
rect -100 -2107 -84 -2073
rect 84 -2107 100 -2073
rect -146 -2157 -112 -2141
rect -146 -2949 -112 -2933
rect 112 -2157 146 -2141
rect 112 -2949 146 -2933
rect -100 -3017 -84 -2983
rect 84 -3017 100 -2983
rect -100 -3125 -84 -3091
rect 84 -3125 100 -3091
rect -146 -3175 -112 -3159
rect -146 -3967 -112 -3951
rect 112 -3175 146 -3159
rect 112 -3967 146 -3951
rect -100 -4035 -84 -4001
rect 84 -4035 100 -4001
rect -100 -4143 -84 -4109
rect 84 -4143 100 -4109
rect -146 -4193 -112 -4177
rect -146 -4985 -112 -4969
rect 112 -4193 146 -4177
rect 112 -4985 146 -4969
rect -100 -5053 -84 -5019
rect 84 -5053 100 -5019
rect -100 -5161 -84 -5127
rect 84 -5161 100 -5127
rect -146 -5211 -112 -5195
rect -146 -6003 -112 -5987
rect 112 -5211 146 -5195
rect 112 -6003 146 -5987
rect -100 -6071 -84 -6037
rect 84 -6071 100 -6037
rect -100 -6179 -84 -6145
rect 84 -6179 100 -6145
rect -146 -6229 -112 -6213
rect -146 -7021 -112 -7005
rect 112 -6229 146 -6213
rect 112 -7021 146 -7005
rect -100 -7089 -84 -7055
rect 84 -7089 100 -7055
rect -100 -7197 -84 -7163
rect 84 -7197 100 -7163
rect -146 -7247 -112 -7231
rect -146 -8039 -112 -8023
rect 112 -7247 146 -7231
rect 112 -8039 146 -8023
rect -100 -8107 -84 -8073
rect 84 -8107 100 -8073
rect -100 -8215 -84 -8181
rect 84 -8215 100 -8181
rect -146 -8265 -112 -8249
rect -146 -9057 -112 -9041
rect 112 -8265 146 -8249
rect 112 -9057 146 -9041
rect -100 -9125 -84 -9091
rect 84 -9125 100 -9091
rect -100 -9233 -84 -9199
rect 84 -9233 100 -9199
rect -146 -9283 -112 -9267
rect -146 -10075 -112 -10059
rect 112 -9283 146 -9267
rect 112 -10075 146 -10059
rect -100 -10143 -84 -10109
rect 84 -10143 100 -10109
rect -280 -10247 -246 -10185
rect 246 -10247 280 -10185
rect -280 -10281 -184 -10247
rect 184 -10281 280 -10247
<< viali >>
rect -84 10109 84 10143
rect -146 9283 -112 10059
rect 112 9283 146 10059
rect -84 9199 84 9233
rect -84 9091 84 9125
rect -146 8265 -112 9041
rect 112 8265 146 9041
rect -84 8181 84 8215
rect -84 8073 84 8107
rect -146 7247 -112 8023
rect 112 7247 146 8023
rect -84 7163 84 7197
rect -84 7055 84 7089
rect -146 6229 -112 7005
rect 112 6229 146 7005
rect -84 6145 84 6179
rect -84 6037 84 6071
rect -146 5211 -112 5987
rect 112 5211 146 5987
rect -84 5127 84 5161
rect -84 5019 84 5053
rect -146 4193 -112 4969
rect 112 4193 146 4969
rect -84 4109 84 4143
rect -84 4001 84 4035
rect -146 3175 -112 3951
rect 112 3175 146 3951
rect -84 3091 84 3125
rect -84 2983 84 3017
rect -146 2157 -112 2933
rect 112 2157 146 2933
rect -84 2073 84 2107
rect -84 1965 84 1999
rect -146 1139 -112 1915
rect 112 1139 146 1915
rect -84 1055 84 1089
rect -84 947 84 981
rect -146 121 -112 897
rect 112 121 146 897
rect -84 37 84 71
rect -84 -71 84 -37
rect -146 -897 -112 -121
rect 112 -897 146 -121
rect -84 -981 84 -947
rect -84 -1089 84 -1055
rect -146 -1915 -112 -1139
rect 112 -1915 146 -1139
rect -84 -1999 84 -1965
rect -84 -2107 84 -2073
rect -146 -2933 -112 -2157
rect 112 -2933 146 -2157
rect -84 -3017 84 -2983
rect -84 -3125 84 -3091
rect -146 -3951 -112 -3175
rect 112 -3951 146 -3175
rect -84 -4035 84 -4001
rect -84 -4143 84 -4109
rect -146 -4969 -112 -4193
rect 112 -4969 146 -4193
rect -84 -5053 84 -5019
rect -84 -5161 84 -5127
rect -146 -5987 -112 -5211
rect 112 -5987 146 -5211
rect -84 -6071 84 -6037
rect -84 -6179 84 -6145
rect -146 -7005 -112 -6229
rect 112 -7005 146 -6229
rect -84 -7089 84 -7055
rect -84 -7197 84 -7163
rect -146 -8023 -112 -7247
rect 112 -8023 146 -7247
rect -84 -8107 84 -8073
rect -84 -8215 84 -8181
rect -146 -9041 -112 -8265
rect 112 -9041 146 -8265
rect -84 -9125 84 -9091
rect -84 -9233 84 -9199
rect -146 -10059 -112 -9283
rect 112 -10059 146 -9283
rect -84 -10143 84 -10109
<< metal1 >>
rect -96 10143 96 10149
rect -96 10109 -84 10143
rect 84 10109 96 10143
rect -96 10103 96 10109
rect -152 10059 -106 10071
rect -152 9283 -146 10059
rect -112 9283 -106 10059
rect -152 9271 -106 9283
rect 106 10059 152 10071
rect 106 9283 112 10059
rect 146 9283 152 10059
rect 106 9271 152 9283
rect -96 9233 96 9239
rect -96 9199 -84 9233
rect 84 9199 96 9233
rect -96 9193 96 9199
rect -96 9125 96 9131
rect -96 9091 -84 9125
rect 84 9091 96 9125
rect -96 9085 96 9091
rect -152 9041 -106 9053
rect -152 8265 -146 9041
rect -112 8265 -106 9041
rect -152 8253 -106 8265
rect 106 9041 152 9053
rect 106 8265 112 9041
rect 146 8265 152 9041
rect 106 8253 152 8265
rect -96 8215 96 8221
rect -96 8181 -84 8215
rect 84 8181 96 8215
rect -96 8175 96 8181
rect -96 8107 96 8113
rect -96 8073 -84 8107
rect 84 8073 96 8107
rect -96 8067 96 8073
rect -152 8023 -106 8035
rect -152 7247 -146 8023
rect -112 7247 -106 8023
rect -152 7235 -106 7247
rect 106 8023 152 8035
rect 106 7247 112 8023
rect 146 7247 152 8023
rect 106 7235 152 7247
rect -96 7197 96 7203
rect -96 7163 -84 7197
rect 84 7163 96 7197
rect -96 7157 96 7163
rect -96 7089 96 7095
rect -96 7055 -84 7089
rect 84 7055 96 7089
rect -96 7049 96 7055
rect -152 7005 -106 7017
rect -152 6229 -146 7005
rect -112 6229 -106 7005
rect -152 6217 -106 6229
rect 106 7005 152 7017
rect 106 6229 112 7005
rect 146 6229 152 7005
rect 106 6217 152 6229
rect -96 6179 96 6185
rect -96 6145 -84 6179
rect 84 6145 96 6179
rect -96 6139 96 6145
rect -96 6071 96 6077
rect -96 6037 -84 6071
rect 84 6037 96 6071
rect -96 6031 96 6037
rect -152 5987 -106 5999
rect -152 5211 -146 5987
rect -112 5211 -106 5987
rect -152 5199 -106 5211
rect 106 5987 152 5999
rect 106 5211 112 5987
rect 146 5211 152 5987
rect 106 5199 152 5211
rect -96 5161 96 5167
rect -96 5127 -84 5161
rect 84 5127 96 5161
rect -96 5121 96 5127
rect -96 5053 96 5059
rect -96 5019 -84 5053
rect 84 5019 96 5053
rect -96 5013 96 5019
rect -152 4969 -106 4981
rect -152 4193 -146 4969
rect -112 4193 -106 4969
rect -152 4181 -106 4193
rect 106 4969 152 4981
rect 106 4193 112 4969
rect 146 4193 152 4969
rect 106 4181 152 4193
rect -96 4143 96 4149
rect -96 4109 -84 4143
rect 84 4109 96 4143
rect -96 4103 96 4109
rect -96 4035 96 4041
rect -96 4001 -84 4035
rect 84 4001 96 4035
rect -96 3995 96 4001
rect -152 3951 -106 3963
rect -152 3175 -146 3951
rect -112 3175 -106 3951
rect -152 3163 -106 3175
rect 106 3951 152 3963
rect 106 3175 112 3951
rect 146 3175 152 3951
rect 106 3163 152 3175
rect -96 3125 96 3131
rect -96 3091 -84 3125
rect 84 3091 96 3125
rect -96 3085 96 3091
rect -96 3017 96 3023
rect -96 2983 -84 3017
rect 84 2983 96 3017
rect -96 2977 96 2983
rect -152 2933 -106 2945
rect -152 2157 -146 2933
rect -112 2157 -106 2933
rect -152 2145 -106 2157
rect 106 2933 152 2945
rect 106 2157 112 2933
rect 146 2157 152 2933
rect 106 2145 152 2157
rect -96 2107 96 2113
rect -96 2073 -84 2107
rect 84 2073 96 2107
rect -96 2067 96 2073
rect -96 1999 96 2005
rect -96 1965 -84 1999
rect 84 1965 96 1999
rect -96 1959 96 1965
rect -152 1915 -106 1927
rect -152 1139 -146 1915
rect -112 1139 -106 1915
rect -152 1127 -106 1139
rect 106 1915 152 1927
rect 106 1139 112 1915
rect 146 1139 152 1915
rect 106 1127 152 1139
rect -96 1089 96 1095
rect -96 1055 -84 1089
rect 84 1055 96 1089
rect -96 1049 96 1055
rect -96 981 96 987
rect -96 947 -84 981
rect 84 947 96 981
rect -96 941 96 947
rect -152 897 -106 909
rect -152 121 -146 897
rect -112 121 -106 897
rect -152 109 -106 121
rect 106 897 152 909
rect 106 121 112 897
rect 146 121 152 897
rect 106 109 152 121
rect -96 71 96 77
rect -96 37 -84 71
rect 84 37 96 71
rect -96 31 96 37
rect -96 -37 96 -31
rect -96 -71 -84 -37
rect 84 -71 96 -37
rect -96 -77 96 -71
rect -152 -121 -106 -109
rect -152 -897 -146 -121
rect -112 -897 -106 -121
rect -152 -909 -106 -897
rect 106 -121 152 -109
rect 106 -897 112 -121
rect 146 -897 152 -121
rect 106 -909 152 -897
rect -96 -947 96 -941
rect -96 -981 -84 -947
rect 84 -981 96 -947
rect -96 -987 96 -981
rect -96 -1055 96 -1049
rect -96 -1089 -84 -1055
rect 84 -1089 96 -1055
rect -96 -1095 96 -1089
rect -152 -1139 -106 -1127
rect -152 -1915 -146 -1139
rect -112 -1915 -106 -1139
rect -152 -1927 -106 -1915
rect 106 -1139 152 -1127
rect 106 -1915 112 -1139
rect 146 -1915 152 -1139
rect 106 -1927 152 -1915
rect -96 -1965 96 -1959
rect -96 -1999 -84 -1965
rect 84 -1999 96 -1965
rect -96 -2005 96 -1999
rect -96 -2073 96 -2067
rect -96 -2107 -84 -2073
rect 84 -2107 96 -2073
rect -96 -2113 96 -2107
rect -152 -2157 -106 -2145
rect -152 -2933 -146 -2157
rect -112 -2933 -106 -2157
rect -152 -2945 -106 -2933
rect 106 -2157 152 -2145
rect 106 -2933 112 -2157
rect 146 -2933 152 -2157
rect 106 -2945 152 -2933
rect -96 -2983 96 -2977
rect -96 -3017 -84 -2983
rect 84 -3017 96 -2983
rect -96 -3023 96 -3017
rect -96 -3091 96 -3085
rect -96 -3125 -84 -3091
rect 84 -3125 96 -3091
rect -96 -3131 96 -3125
rect -152 -3175 -106 -3163
rect -152 -3951 -146 -3175
rect -112 -3951 -106 -3175
rect -152 -3963 -106 -3951
rect 106 -3175 152 -3163
rect 106 -3951 112 -3175
rect 146 -3951 152 -3175
rect 106 -3963 152 -3951
rect -96 -4001 96 -3995
rect -96 -4035 -84 -4001
rect 84 -4035 96 -4001
rect -96 -4041 96 -4035
rect -96 -4109 96 -4103
rect -96 -4143 -84 -4109
rect 84 -4143 96 -4109
rect -96 -4149 96 -4143
rect -152 -4193 -106 -4181
rect -152 -4969 -146 -4193
rect -112 -4969 -106 -4193
rect -152 -4981 -106 -4969
rect 106 -4193 152 -4181
rect 106 -4969 112 -4193
rect 146 -4969 152 -4193
rect 106 -4981 152 -4969
rect -96 -5019 96 -5013
rect -96 -5053 -84 -5019
rect 84 -5053 96 -5019
rect -96 -5059 96 -5053
rect -96 -5127 96 -5121
rect -96 -5161 -84 -5127
rect 84 -5161 96 -5127
rect -96 -5167 96 -5161
rect -152 -5211 -106 -5199
rect -152 -5987 -146 -5211
rect -112 -5987 -106 -5211
rect -152 -5999 -106 -5987
rect 106 -5211 152 -5199
rect 106 -5987 112 -5211
rect 146 -5987 152 -5211
rect 106 -5999 152 -5987
rect -96 -6037 96 -6031
rect -96 -6071 -84 -6037
rect 84 -6071 96 -6037
rect -96 -6077 96 -6071
rect -96 -6145 96 -6139
rect -96 -6179 -84 -6145
rect 84 -6179 96 -6145
rect -96 -6185 96 -6179
rect -152 -6229 -106 -6217
rect -152 -7005 -146 -6229
rect -112 -7005 -106 -6229
rect -152 -7017 -106 -7005
rect 106 -6229 152 -6217
rect 106 -7005 112 -6229
rect 146 -7005 152 -6229
rect 106 -7017 152 -7005
rect -96 -7055 96 -7049
rect -96 -7089 -84 -7055
rect 84 -7089 96 -7055
rect -96 -7095 96 -7089
rect -96 -7163 96 -7157
rect -96 -7197 -84 -7163
rect 84 -7197 96 -7163
rect -96 -7203 96 -7197
rect -152 -7247 -106 -7235
rect -152 -8023 -146 -7247
rect -112 -8023 -106 -7247
rect -152 -8035 -106 -8023
rect 106 -7247 152 -7235
rect 106 -8023 112 -7247
rect 146 -8023 152 -7247
rect 106 -8035 152 -8023
rect -96 -8073 96 -8067
rect -96 -8107 -84 -8073
rect 84 -8107 96 -8073
rect -96 -8113 96 -8107
rect -96 -8181 96 -8175
rect -96 -8215 -84 -8181
rect 84 -8215 96 -8181
rect -96 -8221 96 -8215
rect -152 -8265 -106 -8253
rect -152 -9041 -146 -8265
rect -112 -9041 -106 -8265
rect -152 -9053 -106 -9041
rect 106 -8265 152 -8253
rect 106 -9041 112 -8265
rect 146 -9041 152 -8265
rect 106 -9053 152 -9041
rect -96 -9091 96 -9085
rect -96 -9125 -84 -9091
rect 84 -9125 96 -9091
rect -96 -9131 96 -9125
rect -96 -9199 96 -9193
rect -96 -9233 -84 -9199
rect 84 -9233 96 -9199
rect -96 -9239 96 -9233
rect -152 -9283 -106 -9271
rect -152 -10059 -146 -9283
rect -112 -10059 -106 -9283
rect -152 -10071 -106 -10059
rect 106 -9283 152 -9271
rect 106 -10059 112 -9283
rect 146 -10059 152 -9283
rect 106 -10071 152 -10059
rect -96 -10109 96 -10103
rect -96 -10143 -84 -10109
rect 84 -10143 96 -10109
rect -96 -10149 96 -10143
<< properties >>
string FIXED_BBOX -263 -10264 263 10264
string gencell sky130_fd_pr__nfet_g5v0d10v5
string library sky130
string parameters w 4.0 l 1.0 m 20 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
