magic
tech sky130A
magscale 1 2
timestamp 1716810006
<< locali >>
rect -17 583 17 617
<< metal1 >>
rect 92 784 136 2260
rect 192 714 238 2318
rect 292 786 336 2262
use sky130_fd_pr__nfet_g5v0d10v5_RVEQ2N  XM1
timestamp 1716808352
transform 1 0 213 0 1 1520
box -278 -985 278 985
<< labels >>
rlabel metal1 98 1502 130 1536 0 D
port 1 nsew
rlabel metal1 200 1502 232 1536 0 G
port 2 nsew
rlabel metal1 298 1504 330 1538 0 S
port 3 nsew
rlabel locali -17 583 17 617 0 B
port 4 nsew
<< end >>
