magic
tech sky130A
magscale 1 2
timestamp 1716807968
<< pwell >>
rect -328 -2185 328 2185
<< mvnmos >>
rect -100 1127 100 1927
rect -100 109 100 909
rect -100 -909 100 -109
rect -100 -1927 100 -1127
<< mvndiff >>
rect -158 1915 -100 1927
rect -158 1139 -146 1915
rect -112 1139 -100 1915
rect -158 1127 -100 1139
rect 100 1915 158 1927
rect 100 1139 112 1915
rect 146 1139 158 1915
rect 100 1127 158 1139
rect -158 897 -100 909
rect -158 121 -146 897
rect -112 121 -100 897
rect -158 109 -100 121
rect 100 897 158 909
rect 100 121 112 897
rect 146 121 158 897
rect 100 109 158 121
rect -158 -121 -100 -109
rect -158 -897 -146 -121
rect -112 -897 -100 -121
rect -158 -909 -100 -897
rect 100 -121 158 -109
rect 100 -897 112 -121
rect 146 -897 158 -121
rect 100 -909 158 -897
rect -158 -1139 -100 -1127
rect -158 -1915 -146 -1139
rect -112 -1915 -100 -1139
rect -158 -1927 -100 -1915
rect 100 -1139 158 -1127
rect 100 -1915 112 -1139
rect 146 -1915 158 -1139
rect 100 -1927 158 -1915
<< mvndiffc >>
rect -146 1139 -112 1915
rect 112 1139 146 1915
rect -146 121 -112 897
rect 112 121 146 897
rect -146 -897 -112 -121
rect 112 -897 146 -121
rect -146 -1915 -112 -1139
rect 112 -1915 146 -1139
<< mvpsubdiff >>
rect -292 2137 292 2149
rect -292 2103 -184 2137
rect 184 2103 292 2137
rect -292 2091 292 2103
rect -292 2041 -234 2091
rect -292 -2041 -280 2041
rect -246 -2041 -234 2041
rect 234 2041 292 2091
rect -292 -2091 -234 -2041
rect 234 -2041 246 2041
rect 280 -2041 292 2041
rect 234 -2091 292 -2041
rect -292 -2103 292 -2091
rect -292 -2137 -184 -2103
rect 184 -2137 292 -2103
rect -292 -2149 292 -2137
<< mvpsubdiffcont >>
rect -184 2103 184 2137
rect -280 -2041 -246 2041
rect 246 -2041 280 2041
rect -184 -2137 184 -2103
<< poly >>
rect -100 1999 100 2015
rect -100 1965 -84 1999
rect 84 1965 100 1999
rect -100 1927 100 1965
rect -100 1089 100 1127
rect -100 1055 -84 1089
rect 84 1055 100 1089
rect -100 1039 100 1055
rect -100 981 100 997
rect -100 947 -84 981
rect 84 947 100 981
rect -100 909 100 947
rect -100 71 100 109
rect -100 37 -84 71
rect 84 37 100 71
rect -100 21 100 37
rect -100 -37 100 -21
rect -100 -71 -84 -37
rect 84 -71 100 -37
rect -100 -109 100 -71
rect -100 -947 100 -909
rect -100 -981 -84 -947
rect 84 -981 100 -947
rect -100 -997 100 -981
rect -100 -1055 100 -1039
rect -100 -1089 -84 -1055
rect 84 -1089 100 -1055
rect -100 -1127 100 -1089
rect -100 -1965 100 -1927
rect -100 -1999 -84 -1965
rect 84 -1999 100 -1965
rect -100 -2015 100 -1999
<< polycont >>
rect -84 1965 84 1999
rect -84 1055 84 1089
rect -84 947 84 981
rect -84 37 84 71
rect -84 -71 84 -37
rect -84 -981 84 -947
rect -84 -1089 84 -1055
rect -84 -1999 84 -1965
<< locali >>
rect -280 2103 -184 2137
rect 184 2103 280 2137
rect -280 2041 -246 2103
rect 246 2041 280 2103
rect -100 1965 -84 1999
rect 84 1965 100 1999
rect -146 1915 -112 1931
rect -146 1123 -112 1139
rect 112 1915 146 1931
rect 112 1123 146 1139
rect -100 1055 -84 1089
rect 84 1055 100 1089
rect -100 947 -84 981
rect 84 947 100 981
rect -146 897 -112 913
rect -146 105 -112 121
rect 112 897 146 913
rect 112 105 146 121
rect -100 37 -84 71
rect 84 37 100 71
rect -100 -71 -84 -37
rect 84 -71 100 -37
rect -146 -121 -112 -105
rect -146 -913 -112 -897
rect 112 -121 146 -105
rect 112 -913 146 -897
rect -100 -981 -84 -947
rect 84 -981 100 -947
rect -100 -1089 -84 -1055
rect 84 -1089 100 -1055
rect -146 -1139 -112 -1123
rect -146 -1931 -112 -1915
rect 112 -1139 146 -1123
rect 112 -1931 146 -1915
rect -100 -1999 -84 -1965
rect 84 -1999 100 -1965
rect -280 -2103 -246 -2041
rect 246 -2103 280 -2041
rect -280 -2137 -184 -2103
rect 184 -2137 280 -2103
<< viali >>
rect -84 1965 84 1999
rect -146 1139 -112 1915
rect 112 1139 146 1915
rect -84 1055 84 1089
rect -84 947 84 981
rect -146 121 -112 897
rect 112 121 146 897
rect -84 37 84 71
rect -84 -71 84 -37
rect -146 -897 -112 -121
rect 112 -897 146 -121
rect -84 -981 84 -947
rect -84 -1089 84 -1055
rect -146 -1915 -112 -1139
rect 112 -1915 146 -1139
rect -84 -1999 84 -1965
<< metal1 >>
rect -96 1999 96 2005
rect -96 1965 -84 1999
rect 84 1965 96 1999
rect -96 1959 96 1965
rect -152 1915 -106 1927
rect -152 1139 -146 1915
rect -112 1139 -106 1915
rect -152 1127 -106 1139
rect 106 1915 152 1927
rect 106 1139 112 1915
rect 146 1139 152 1915
rect 106 1127 152 1139
rect -96 1089 96 1095
rect -96 1055 -84 1089
rect 84 1055 96 1089
rect -96 1049 96 1055
rect -96 981 96 987
rect -96 947 -84 981
rect 84 947 96 981
rect -96 941 96 947
rect -152 897 -106 909
rect -152 121 -146 897
rect -112 121 -106 897
rect -152 109 -106 121
rect 106 897 152 909
rect 106 121 112 897
rect 146 121 152 897
rect 106 109 152 121
rect -96 71 96 77
rect -96 37 -84 71
rect 84 37 96 71
rect -96 31 96 37
rect -96 -37 96 -31
rect -96 -71 -84 -37
rect 84 -71 96 -37
rect -96 -77 96 -71
rect -152 -121 -106 -109
rect -152 -897 -146 -121
rect -112 -897 -106 -121
rect -152 -909 -106 -897
rect 106 -121 152 -109
rect 106 -897 112 -121
rect 146 -897 152 -121
rect 106 -909 152 -897
rect -96 -947 96 -941
rect -96 -981 -84 -947
rect 84 -981 96 -947
rect -96 -987 96 -981
rect -96 -1055 96 -1049
rect -96 -1089 -84 -1055
rect 84 -1089 96 -1055
rect -96 -1095 96 -1089
rect -152 -1139 -106 -1127
rect -152 -1915 -146 -1139
rect -112 -1915 -106 -1139
rect -152 -1927 -106 -1915
rect 106 -1139 152 -1127
rect 106 -1915 112 -1139
rect 146 -1915 152 -1139
rect 106 -1927 152 -1915
rect -96 -1965 96 -1959
rect -96 -1999 -84 -1965
rect 84 -1999 96 -1965
rect -96 -2005 96 -1999
<< properties >>
string FIXED_BBOX -263 -2120 263 2120
string gencell sky130_fd_pr__nfet_g5v0d10v5
string library sky130
string parameters w 4.0 l 1.0 m 4 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
