magic
tech sky130A
magscale 1 2
timestamp 1717127688
<< nwell >>
rect -487 -1762 487 1762
<< mvpmos >>
rect -229 -1536 -29 1464
rect 29 -1536 229 1464
<< mvpdiff >>
rect -287 1452 -229 1464
rect -287 -1524 -275 1452
rect -241 -1524 -229 1452
rect -287 -1536 -229 -1524
rect -29 1452 29 1464
rect -29 -1524 -17 1452
rect 17 -1524 29 1452
rect -29 -1536 29 -1524
rect 229 1452 287 1464
rect 229 -1524 241 1452
rect 275 -1524 287 1452
rect 229 -1536 287 -1524
<< mvpdiffc >>
rect -275 -1524 -241 1452
rect -17 -1524 17 1452
rect 241 -1524 275 1452
<< mvnsubdiff >>
rect -421 1684 421 1696
rect -421 1650 -313 1684
rect 313 1650 421 1684
rect -421 1638 421 1650
rect -421 1588 -363 1638
rect -421 -1588 -409 1588
rect -375 -1588 -363 1588
rect 363 1588 421 1638
rect -421 -1638 -363 -1588
rect 363 -1588 375 1588
rect 409 -1588 421 1588
rect 363 -1638 421 -1588
rect -421 -1650 421 -1638
rect -421 -1684 -313 -1650
rect 313 -1684 421 -1650
rect -421 -1696 421 -1684
<< mvnsubdiffcont >>
rect -313 1650 313 1684
rect -409 -1588 -375 1588
rect 375 -1588 409 1588
rect -313 -1684 313 -1650
<< poly >>
rect -229 1545 -29 1561
rect -229 1511 -213 1545
rect -45 1511 -29 1545
rect -229 1464 -29 1511
rect 29 1545 229 1561
rect 29 1511 45 1545
rect 213 1511 229 1545
rect 29 1464 229 1511
rect -229 -1562 -29 -1536
rect 29 -1562 229 -1536
<< polycont >>
rect -213 1511 -45 1545
rect 45 1511 213 1545
<< locali >>
rect -409 1650 -313 1684
rect 313 1650 409 1684
rect -409 1588 -375 1650
rect 375 1588 409 1650
rect -229 1511 -213 1545
rect -45 1511 -29 1545
rect 29 1511 45 1545
rect 213 1511 229 1545
rect -275 1452 -241 1468
rect -275 -1540 -241 -1524
rect -17 1452 17 1468
rect -17 -1540 17 -1524
rect 241 1452 275 1468
rect 241 -1540 275 -1524
rect -409 -1650 -375 -1588
rect 375 -1650 409 -1588
rect -409 -1684 -313 -1650
rect 313 -1684 409 -1650
<< viali >>
rect -213 1511 -45 1545
rect 45 1511 213 1545
rect -275 -1524 -241 1452
rect -17 -1524 17 1452
rect 241 -1524 275 1452
<< metal1 >>
rect -225 1545 -33 1551
rect -225 1511 -213 1545
rect -45 1511 -33 1545
rect -225 1505 -33 1511
rect 33 1545 225 1551
rect 33 1511 45 1545
rect 213 1511 225 1545
rect 33 1505 225 1511
rect -281 1452 -235 1464
rect -281 -1524 -275 1452
rect -241 -1524 -235 1452
rect -281 -1536 -235 -1524
rect -23 1452 23 1464
rect -23 -1524 -17 1452
rect 17 -1524 23 1452
rect -23 -1536 23 -1524
rect 235 1452 281 1464
rect 235 -1524 241 1452
rect 275 -1524 281 1452
rect 235 -1536 281 -1524
<< properties >>
string FIXED_BBOX -392 -1667 392 1667
string gencell sky130_fd_pr__pfet_g5v0d10v5
string library sky130
string parameters w 15.0 l 1.0 m 1 nf 2 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
