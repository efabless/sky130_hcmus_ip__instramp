magic
tech sky130A
magscale 1 2
timestamp 1716807968
<< pwell >>
rect -328 -4221 328 4221
<< mvnmos >>
rect -100 3163 100 3963
rect -100 2145 100 2945
rect -100 1127 100 1927
rect -100 109 100 909
rect -100 -909 100 -109
rect -100 -1927 100 -1127
rect -100 -2945 100 -2145
rect -100 -3963 100 -3163
<< mvndiff >>
rect -158 3951 -100 3963
rect -158 3175 -146 3951
rect -112 3175 -100 3951
rect -158 3163 -100 3175
rect 100 3951 158 3963
rect 100 3175 112 3951
rect 146 3175 158 3951
rect 100 3163 158 3175
rect -158 2933 -100 2945
rect -158 2157 -146 2933
rect -112 2157 -100 2933
rect -158 2145 -100 2157
rect 100 2933 158 2945
rect 100 2157 112 2933
rect 146 2157 158 2933
rect 100 2145 158 2157
rect -158 1915 -100 1927
rect -158 1139 -146 1915
rect -112 1139 -100 1915
rect -158 1127 -100 1139
rect 100 1915 158 1927
rect 100 1139 112 1915
rect 146 1139 158 1915
rect 100 1127 158 1139
rect -158 897 -100 909
rect -158 121 -146 897
rect -112 121 -100 897
rect -158 109 -100 121
rect 100 897 158 909
rect 100 121 112 897
rect 146 121 158 897
rect 100 109 158 121
rect -158 -121 -100 -109
rect -158 -897 -146 -121
rect -112 -897 -100 -121
rect -158 -909 -100 -897
rect 100 -121 158 -109
rect 100 -897 112 -121
rect 146 -897 158 -121
rect 100 -909 158 -897
rect -158 -1139 -100 -1127
rect -158 -1915 -146 -1139
rect -112 -1915 -100 -1139
rect -158 -1927 -100 -1915
rect 100 -1139 158 -1127
rect 100 -1915 112 -1139
rect 146 -1915 158 -1139
rect 100 -1927 158 -1915
rect -158 -2157 -100 -2145
rect -158 -2933 -146 -2157
rect -112 -2933 -100 -2157
rect -158 -2945 -100 -2933
rect 100 -2157 158 -2145
rect 100 -2933 112 -2157
rect 146 -2933 158 -2157
rect 100 -2945 158 -2933
rect -158 -3175 -100 -3163
rect -158 -3951 -146 -3175
rect -112 -3951 -100 -3175
rect -158 -3963 -100 -3951
rect 100 -3175 158 -3163
rect 100 -3951 112 -3175
rect 146 -3951 158 -3175
rect 100 -3963 158 -3951
<< mvndiffc >>
rect -146 3175 -112 3951
rect 112 3175 146 3951
rect -146 2157 -112 2933
rect 112 2157 146 2933
rect -146 1139 -112 1915
rect 112 1139 146 1915
rect -146 121 -112 897
rect 112 121 146 897
rect -146 -897 -112 -121
rect 112 -897 146 -121
rect -146 -1915 -112 -1139
rect 112 -1915 146 -1139
rect -146 -2933 -112 -2157
rect 112 -2933 146 -2157
rect -146 -3951 -112 -3175
rect 112 -3951 146 -3175
<< mvpsubdiff >>
rect -292 4173 292 4185
rect -292 4139 -184 4173
rect 184 4139 292 4173
rect -292 4127 292 4139
rect -292 4077 -234 4127
rect -292 -4077 -280 4077
rect -246 -4077 -234 4077
rect 234 4077 292 4127
rect -292 -4127 -234 -4077
rect 234 -4077 246 4077
rect 280 -4077 292 4077
rect 234 -4127 292 -4077
rect -292 -4139 292 -4127
rect -292 -4173 -184 -4139
rect 184 -4173 292 -4139
rect -292 -4185 292 -4173
<< mvpsubdiffcont >>
rect -184 4139 184 4173
rect -280 -4077 -246 4077
rect 246 -4077 280 4077
rect -184 -4173 184 -4139
<< poly >>
rect -100 4035 100 4051
rect -100 4001 -84 4035
rect 84 4001 100 4035
rect -100 3963 100 4001
rect -100 3125 100 3163
rect -100 3091 -84 3125
rect 84 3091 100 3125
rect -100 3075 100 3091
rect -100 3017 100 3033
rect -100 2983 -84 3017
rect 84 2983 100 3017
rect -100 2945 100 2983
rect -100 2107 100 2145
rect -100 2073 -84 2107
rect 84 2073 100 2107
rect -100 2057 100 2073
rect -100 1999 100 2015
rect -100 1965 -84 1999
rect 84 1965 100 1999
rect -100 1927 100 1965
rect -100 1089 100 1127
rect -100 1055 -84 1089
rect 84 1055 100 1089
rect -100 1039 100 1055
rect -100 981 100 997
rect -100 947 -84 981
rect 84 947 100 981
rect -100 909 100 947
rect -100 71 100 109
rect -100 37 -84 71
rect 84 37 100 71
rect -100 21 100 37
rect -100 -37 100 -21
rect -100 -71 -84 -37
rect 84 -71 100 -37
rect -100 -109 100 -71
rect -100 -947 100 -909
rect -100 -981 -84 -947
rect 84 -981 100 -947
rect -100 -997 100 -981
rect -100 -1055 100 -1039
rect -100 -1089 -84 -1055
rect 84 -1089 100 -1055
rect -100 -1127 100 -1089
rect -100 -1965 100 -1927
rect -100 -1999 -84 -1965
rect 84 -1999 100 -1965
rect -100 -2015 100 -1999
rect -100 -2073 100 -2057
rect -100 -2107 -84 -2073
rect 84 -2107 100 -2073
rect -100 -2145 100 -2107
rect -100 -2983 100 -2945
rect -100 -3017 -84 -2983
rect 84 -3017 100 -2983
rect -100 -3033 100 -3017
rect -100 -3091 100 -3075
rect -100 -3125 -84 -3091
rect 84 -3125 100 -3091
rect -100 -3163 100 -3125
rect -100 -4001 100 -3963
rect -100 -4035 -84 -4001
rect 84 -4035 100 -4001
rect -100 -4051 100 -4035
<< polycont >>
rect -84 4001 84 4035
rect -84 3091 84 3125
rect -84 2983 84 3017
rect -84 2073 84 2107
rect -84 1965 84 1999
rect -84 1055 84 1089
rect -84 947 84 981
rect -84 37 84 71
rect -84 -71 84 -37
rect -84 -981 84 -947
rect -84 -1089 84 -1055
rect -84 -1999 84 -1965
rect -84 -2107 84 -2073
rect -84 -3017 84 -2983
rect -84 -3125 84 -3091
rect -84 -4035 84 -4001
<< locali >>
rect -280 4139 -184 4173
rect 184 4139 280 4173
rect -280 4077 -246 4139
rect 246 4077 280 4139
rect -100 4001 -84 4035
rect 84 4001 100 4035
rect -146 3951 -112 3967
rect -146 3159 -112 3175
rect 112 3951 146 3967
rect 112 3159 146 3175
rect -100 3091 -84 3125
rect 84 3091 100 3125
rect -100 2983 -84 3017
rect 84 2983 100 3017
rect -146 2933 -112 2949
rect -146 2141 -112 2157
rect 112 2933 146 2949
rect 112 2141 146 2157
rect -100 2073 -84 2107
rect 84 2073 100 2107
rect -100 1965 -84 1999
rect 84 1965 100 1999
rect -146 1915 -112 1931
rect -146 1123 -112 1139
rect 112 1915 146 1931
rect 112 1123 146 1139
rect -100 1055 -84 1089
rect 84 1055 100 1089
rect -100 947 -84 981
rect 84 947 100 981
rect -146 897 -112 913
rect -146 105 -112 121
rect 112 897 146 913
rect 112 105 146 121
rect -100 37 -84 71
rect 84 37 100 71
rect -100 -71 -84 -37
rect 84 -71 100 -37
rect -146 -121 -112 -105
rect -146 -913 -112 -897
rect 112 -121 146 -105
rect 112 -913 146 -897
rect -100 -981 -84 -947
rect 84 -981 100 -947
rect -100 -1089 -84 -1055
rect 84 -1089 100 -1055
rect -146 -1139 -112 -1123
rect -146 -1931 -112 -1915
rect 112 -1139 146 -1123
rect 112 -1931 146 -1915
rect -100 -1999 -84 -1965
rect 84 -1999 100 -1965
rect -100 -2107 -84 -2073
rect 84 -2107 100 -2073
rect -146 -2157 -112 -2141
rect -146 -2949 -112 -2933
rect 112 -2157 146 -2141
rect 112 -2949 146 -2933
rect -100 -3017 -84 -2983
rect 84 -3017 100 -2983
rect -100 -3125 -84 -3091
rect 84 -3125 100 -3091
rect -146 -3175 -112 -3159
rect -146 -3967 -112 -3951
rect 112 -3175 146 -3159
rect 112 -3967 146 -3951
rect -100 -4035 -84 -4001
rect 84 -4035 100 -4001
rect -280 -4139 -246 -4077
rect 246 -4139 280 -4077
rect -280 -4173 -184 -4139
rect 184 -4173 280 -4139
<< viali >>
rect -84 4001 84 4035
rect -146 3175 -112 3951
rect 112 3175 146 3951
rect -84 3091 84 3125
rect -84 2983 84 3017
rect -146 2157 -112 2933
rect 112 2157 146 2933
rect -84 2073 84 2107
rect -84 1965 84 1999
rect -146 1139 -112 1915
rect 112 1139 146 1915
rect -84 1055 84 1089
rect -84 947 84 981
rect -146 121 -112 897
rect 112 121 146 897
rect -84 37 84 71
rect -84 -71 84 -37
rect -146 -897 -112 -121
rect 112 -897 146 -121
rect -84 -981 84 -947
rect -84 -1089 84 -1055
rect -146 -1915 -112 -1139
rect 112 -1915 146 -1139
rect -84 -1999 84 -1965
rect -84 -2107 84 -2073
rect -146 -2933 -112 -2157
rect 112 -2933 146 -2157
rect -84 -3017 84 -2983
rect -84 -3125 84 -3091
rect -146 -3951 -112 -3175
rect 112 -3951 146 -3175
rect -84 -4035 84 -4001
<< metal1 >>
rect -96 4035 96 4041
rect -96 4001 -84 4035
rect 84 4001 96 4035
rect -96 3995 96 4001
rect -152 3951 -106 3963
rect -152 3175 -146 3951
rect -112 3175 -106 3951
rect -152 3163 -106 3175
rect 106 3951 152 3963
rect 106 3175 112 3951
rect 146 3175 152 3951
rect 106 3163 152 3175
rect -96 3125 96 3131
rect -96 3091 -84 3125
rect 84 3091 96 3125
rect -96 3085 96 3091
rect -96 3017 96 3023
rect -96 2983 -84 3017
rect 84 2983 96 3017
rect -96 2977 96 2983
rect -152 2933 -106 2945
rect -152 2157 -146 2933
rect -112 2157 -106 2933
rect -152 2145 -106 2157
rect 106 2933 152 2945
rect 106 2157 112 2933
rect 146 2157 152 2933
rect 106 2145 152 2157
rect -96 2107 96 2113
rect -96 2073 -84 2107
rect 84 2073 96 2107
rect -96 2067 96 2073
rect -96 1999 96 2005
rect -96 1965 -84 1999
rect 84 1965 96 1999
rect -96 1959 96 1965
rect -152 1915 -106 1927
rect -152 1139 -146 1915
rect -112 1139 -106 1915
rect -152 1127 -106 1139
rect 106 1915 152 1927
rect 106 1139 112 1915
rect 146 1139 152 1915
rect 106 1127 152 1139
rect -96 1089 96 1095
rect -96 1055 -84 1089
rect 84 1055 96 1089
rect -96 1049 96 1055
rect -96 981 96 987
rect -96 947 -84 981
rect 84 947 96 981
rect -96 941 96 947
rect -152 897 -106 909
rect -152 121 -146 897
rect -112 121 -106 897
rect -152 109 -106 121
rect 106 897 152 909
rect 106 121 112 897
rect 146 121 152 897
rect 106 109 152 121
rect -96 71 96 77
rect -96 37 -84 71
rect 84 37 96 71
rect -96 31 96 37
rect -96 -37 96 -31
rect -96 -71 -84 -37
rect 84 -71 96 -37
rect -96 -77 96 -71
rect -152 -121 -106 -109
rect -152 -897 -146 -121
rect -112 -897 -106 -121
rect -152 -909 -106 -897
rect 106 -121 152 -109
rect 106 -897 112 -121
rect 146 -897 152 -121
rect 106 -909 152 -897
rect -96 -947 96 -941
rect -96 -981 -84 -947
rect 84 -981 96 -947
rect -96 -987 96 -981
rect -96 -1055 96 -1049
rect -96 -1089 -84 -1055
rect 84 -1089 96 -1055
rect -96 -1095 96 -1089
rect -152 -1139 -106 -1127
rect -152 -1915 -146 -1139
rect -112 -1915 -106 -1139
rect -152 -1927 -106 -1915
rect 106 -1139 152 -1127
rect 106 -1915 112 -1139
rect 146 -1915 152 -1139
rect 106 -1927 152 -1915
rect -96 -1965 96 -1959
rect -96 -1999 -84 -1965
rect 84 -1999 96 -1965
rect -96 -2005 96 -1999
rect -96 -2073 96 -2067
rect -96 -2107 -84 -2073
rect 84 -2107 96 -2073
rect -96 -2113 96 -2107
rect -152 -2157 -106 -2145
rect -152 -2933 -146 -2157
rect -112 -2933 -106 -2157
rect -152 -2945 -106 -2933
rect 106 -2157 152 -2145
rect 106 -2933 112 -2157
rect 146 -2933 152 -2157
rect 106 -2945 152 -2933
rect -96 -2983 96 -2977
rect -96 -3017 -84 -2983
rect 84 -3017 96 -2983
rect -96 -3023 96 -3017
rect -96 -3091 96 -3085
rect -96 -3125 -84 -3091
rect 84 -3125 96 -3091
rect -96 -3131 96 -3125
rect -152 -3175 -106 -3163
rect -152 -3951 -146 -3175
rect -112 -3951 -106 -3175
rect -152 -3963 -106 -3951
rect 106 -3175 152 -3163
rect 106 -3951 112 -3175
rect 146 -3951 152 -3175
rect 106 -3963 152 -3951
rect -96 -4001 96 -3995
rect -96 -4035 -84 -4001
rect 84 -4035 96 -4001
rect -96 -4041 96 -4035
<< properties >>
string FIXED_BBOX -263 -4156 263 4156
string gencell sky130_fd_pr__nfet_g5v0d10v5
string library sky130
string parameters w 4.0 l 1.0 m 8 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
