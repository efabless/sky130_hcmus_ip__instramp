magic
tech sky130A
timestamp 1716175101
<< nmos >>
rect 0 0 15 100
<< ndiff >>
rect -45 85 0 100
rect -45 15 -35 85
rect -15 15 0 85
rect -45 0 0 15
rect 15 85 60 100
rect 15 15 30 85
rect 50 15 60 85
rect 15 0 60 15
<< ndiffc >>
rect -35 15 -15 85
rect 30 15 50 85
<< psubdiff >>
rect -85 85 -45 100
rect -85 15 -75 85
rect -55 15 -45 85
rect -85 0 -45 15
<< psubdiffcont >>
rect -75 15 -55 85
<< poly >>
rect 0 100 15 115
rect 0 -15 15 0
<< locali >>
rect -85 85 -5 90
rect -85 15 -75 85
rect -55 15 -35 85
rect -15 15 -5 85
rect -85 10 -5 15
rect 20 85 60 90
rect 20 15 30 85
rect 50 15 60 85
rect 20 10 60 15
rect -85 5 -35 10
<< end >>
