magic
tech sky130A
magscale 1 2
timestamp 1718246682
<< pwell >>
rect -235 -902 235 902
<< psubdiff >>
rect -199 832 -103 866
rect 103 832 199 866
rect -199 770 -165 832
rect 165 770 199 832
rect -199 -832 -165 -770
rect 165 -832 199 -770
rect -199 -866 -103 -832
rect 103 -866 199 -832
<< psubdiffcont >>
rect -103 832 103 866
rect -199 -770 -165 770
rect 165 -770 199 770
rect -103 -866 103 -832
<< xpolycontact >>
rect -69 304 69 736
rect -69 -736 69 -304
<< ppolyres >>
rect -69 -304 69 304
<< locali >>
rect -199 832 -103 866
rect 103 832 199 866
rect -199 770 -165 832
rect 165 770 199 832
rect -199 -832 -165 -770
rect 165 -832 199 -770
rect -199 -866 -103 -832
rect 103 -866 199 -832
<< viali >>
rect -53 321 53 718
rect -53 -718 53 -321
<< metal1 >>
rect -59 718 59 730
rect -59 321 -53 718
rect 53 321 59 718
rect -59 309 59 321
rect -59 -321 59 -309
rect -59 -718 -53 -321
rect 53 -718 59 -321
rect -59 -730 59 -718
<< properties >>
string FIXED_BBOX -182 -849 182 849
string gencell sky130_fd_pr__res_high_po_0p69
string library sky130
string parameters w 0.69 l 3.20 m 1 nx 1 wmin 0.690 lmin 0.50 rho 319.8 val 2.047k dummy 0 dw 0.0 term 194.82 sterm 0.0 caplen 0 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_high_po_0p35  sky130_fd_pr__res_high_po_0p69 sky130_fd_pr__res_high_po_1p41  sky130_fd_pr__res_high_po_2p85 sky130_fd_pr__res_high_po_5p73} snake 0 full_metal 1 wmax 0.690 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
