magic
tech sky130A
magscale 1 2
timestamp 1720214482
<< nwell >>
rect -487 -397 487 397
<< mvpmos >>
rect -229 -100 -29 100
rect 29 -100 229 100
<< mvpdiff >>
rect -287 88 -229 100
rect -287 -88 -275 88
rect -241 -88 -229 88
rect -287 -100 -229 -88
rect -29 88 29 100
rect -29 -88 -17 88
rect 17 -88 29 88
rect -29 -100 29 -88
rect 229 88 287 100
rect 229 -88 241 88
rect 275 -88 287 88
rect 229 -100 287 -88
<< mvpdiffc >>
rect -275 -88 -241 88
rect -17 -88 17 88
rect 241 -88 275 88
<< mvnsubdiff >>
rect -421 319 421 331
rect -421 285 -313 319
rect 313 285 421 319
rect -421 273 421 285
rect -421 223 -363 273
rect -421 -223 -409 223
rect -375 -223 -363 223
rect 363 223 421 273
rect -421 -273 -363 -223
rect 363 -223 375 223
rect 409 -223 421 223
rect 363 -273 421 -223
rect -421 -285 421 -273
rect -421 -319 -313 -285
rect 313 -319 421 -285
rect -421 -331 421 -319
<< mvnsubdiffcont >>
rect -313 285 313 319
rect -409 -223 -375 223
rect 375 -223 409 223
rect -313 -319 313 -285
<< poly >>
rect -229 181 -29 197
rect -229 147 -213 181
rect -45 147 -29 181
rect -229 100 -29 147
rect 29 181 229 197
rect 29 147 45 181
rect 213 147 229 181
rect 29 100 229 147
rect -229 -147 -29 -100
rect -229 -181 -213 -147
rect -45 -181 -29 -147
rect -229 -197 -29 -181
rect 29 -147 229 -100
rect 29 -181 45 -147
rect 213 -181 229 -147
rect 29 -197 229 -181
<< polycont >>
rect -213 147 -45 181
rect 45 147 213 181
rect -213 -181 -45 -147
rect 45 -181 213 -147
<< locali >>
rect -409 285 -313 319
rect 313 285 409 319
rect -409 223 -375 285
rect 375 223 409 285
rect -229 147 -213 181
rect -45 147 -29 181
rect 29 147 45 181
rect 213 147 229 181
rect -275 88 -241 104
rect -275 -104 -241 -88
rect -17 88 17 104
rect -17 -104 17 -88
rect 241 88 275 104
rect 241 -104 275 -88
rect -229 -181 -213 -147
rect -45 -181 -29 -147
rect 29 -181 45 -147
rect 213 -181 229 -147
rect -409 -285 -375 -223
rect 375 -285 409 -223
rect -409 -319 -313 -285
rect 313 -319 409 -285
<< viali >>
rect -213 147 -45 181
rect 45 147 213 181
rect -275 -88 -241 88
rect -17 -88 17 88
rect 241 -88 275 88
rect -213 -181 -45 -147
rect 45 -181 213 -147
<< metal1 >>
rect -225 181 -33 187
rect -225 147 -213 181
rect -45 147 -33 181
rect -225 141 -33 147
rect 33 181 225 187
rect 33 147 45 181
rect 213 147 225 181
rect 33 141 225 147
rect -281 88 -235 100
rect -281 -88 -275 88
rect -241 -88 -235 88
rect -281 -100 -235 -88
rect -23 88 23 100
rect -23 -88 -17 88
rect 17 -88 23 88
rect -23 -100 23 -88
rect 235 88 281 100
rect 235 -88 241 88
rect 275 -88 281 88
rect 235 -100 281 -88
rect -225 -147 -33 -141
rect -225 -181 -213 -147
rect -45 -181 -33 -147
rect -225 -187 -33 -181
rect 33 -147 225 -141
rect 33 -181 45 -147
rect 213 -181 225 -147
rect 33 -187 225 -181
<< properties >>
string FIXED_BBOX -392 -302 392 302
string gencell sky130_fd_pr__pfet_g5v0d10v5
string library sky130
string parameters w 1 l 1 m 1 nf 2 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
