magic
tech sky130A
magscale 1 2
timestamp 1717127688
<< pwell >>
rect -715 -723 715 723
<< mvnmos >>
rect -487 -465 -287 465
rect -229 -465 -29 465
rect 29 -465 229 465
rect 287 -465 487 465
<< mvndiff >>
rect -545 453 -487 465
rect -545 -453 -533 453
rect -499 -453 -487 453
rect -545 -465 -487 -453
rect -287 453 -229 465
rect -287 -453 -275 453
rect -241 -453 -229 453
rect -287 -465 -229 -453
rect -29 453 29 465
rect -29 -453 -17 453
rect 17 -453 29 453
rect -29 -465 29 -453
rect 229 453 287 465
rect 229 -453 241 453
rect 275 -453 287 453
rect 229 -465 287 -453
rect 487 453 545 465
rect 487 -453 499 453
rect 533 -453 545 453
rect 487 -465 545 -453
<< mvndiffc >>
rect -533 -453 -499 453
rect -275 -453 -241 453
rect -17 -453 17 453
rect 241 -453 275 453
rect 499 -453 533 453
<< mvpsubdiff >>
rect -679 675 679 687
rect -679 641 -571 675
rect 571 641 679 675
rect -679 629 679 641
rect -679 579 -621 629
rect -679 -579 -667 579
rect -633 -579 -621 579
rect 621 579 679 629
rect -679 -629 -621 -579
rect 621 -579 633 579
rect 667 -579 679 579
rect 621 -629 679 -579
rect -679 -641 679 -629
rect -679 -675 -571 -641
rect 571 -675 679 -641
rect -679 -687 679 -675
<< mvpsubdiffcont >>
rect -571 641 571 675
rect -667 -579 -633 579
rect 633 -579 667 579
rect -571 -675 571 -641
<< poly >>
rect -487 537 -287 553
rect -487 503 -471 537
rect -303 503 -287 537
rect -487 465 -287 503
rect -229 537 -29 553
rect -229 503 -213 537
rect -45 503 -29 537
rect -229 465 -29 503
rect 29 537 229 553
rect 29 503 45 537
rect 213 503 229 537
rect 29 465 229 503
rect 287 537 487 553
rect 287 503 303 537
rect 471 503 487 537
rect 287 465 487 503
rect -487 -503 -287 -465
rect -487 -537 -471 -503
rect -303 -537 -287 -503
rect -487 -553 -287 -537
rect -229 -503 -29 -465
rect -229 -537 -213 -503
rect -45 -537 -29 -503
rect -229 -553 -29 -537
rect 29 -503 229 -465
rect 29 -537 45 -503
rect 213 -537 229 -503
rect 29 -553 229 -537
rect 287 -503 487 -465
rect 287 -537 303 -503
rect 471 -537 487 -503
rect 287 -553 487 -537
<< polycont >>
rect -471 503 -303 537
rect -213 503 -45 537
rect 45 503 213 537
rect 303 503 471 537
rect -471 -537 -303 -503
rect -213 -537 -45 -503
rect 45 -537 213 -503
rect 303 -537 471 -503
<< locali >>
rect -667 641 -571 675
rect 571 641 667 675
rect -667 579 -633 641
rect 633 579 667 641
rect -487 503 -471 537
rect -303 503 -287 537
rect -229 503 -213 537
rect -45 503 -29 537
rect 29 503 45 537
rect 213 503 229 537
rect 287 503 303 537
rect 471 503 487 537
rect -533 453 -499 469
rect -533 -469 -499 -453
rect -275 453 -241 469
rect -275 -469 -241 -453
rect -17 453 17 469
rect -17 -469 17 -453
rect 241 453 275 469
rect 241 -469 275 -453
rect 499 453 533 469
rect 499 -469 533 -453
rect -487 -537 -471 -503
rect -303 -537 -287 -503
rect -229 -537 -213 -503
rect -45 -537 -29 -503
rect 29 -537 45 -503
rect 213 -537 229 -503
rect 287 -537 303 -503
rect 471 -537 487 -503
rect -667 -641 -633 -579
rect 633 -641 667 -579
rect -667 -675 -571 -641
rect 571 -675 667 -641
<< viali >>
rect -471 503 -303 537
rect -213 503 -45 537
rect 45 503 213 537
rect 303 503 471 537
rect -533 -453 -499 453
rect -275 -453 -241 453
rect -17 -453 17 453
rect 241 -453 275 453
rect 499 -453 533 453
rect -471 -537 -303 -503
rect -213 -537 -45 -503
rect 45 -537 213 -503
rect 303 -537 471 -503
<< metal1 >>
rect -483 537 -291 543
rect -483 503 -471 537
rect -303 503 -291 537
rect -483 497 -291 503
rect -225 537 -33 543
rect -225 503 -213 537
rect -45 503 -33 537
rect -225 497 -33 503
rect 33 537 225 543
rect 33 503 45 537
rect 213 503 225 537
rect 33 497 225 503
rect 291 537 483 543
rect 291 503 303 537
rect 471 503 483 537
rect 291 497 483 503
rect -539 453 -493 465
rect -539 -453 -533 453
rect -499 -453 -493 453
rect -539 -465 -493 -453
rect -281 453 -235 465
rect -281 -453 -275 453
rect -241 -453 -235 453
rect -281 -465 -235 -453
rect -23 453 23 465
rect -23 -453 -17 453
rect 17 -453 23 453
rect -23 -465 23 -453
rect 235 453 281 465
rect 235 -453 241 453
rect 275 -453 281 453
rect 235 -465 281 -453
rect 493 453 539 465
rect 493 -453 499 453
rect 533 -453 539 453
rect 493 -465 539 -453
rect -483 -503 -291 -497
rect -483 -537 -471 -503
rect -303 -537 -291 -503
rect -483 -543 -291 -537
rect -225 -503 -33 -497
rect -225 -537 -213 -503
rect -45 -537 -33 -503
rect -225 -543 -33 -537
rect 33 -503 225 -497
rect 33 -537 45 -503
rect 213 -537 225 -503
rect 33 -543 225 -537
rect 291 -503 483 -497
rect 291 -537 303 -503
rect 471 -537 483 -503
rect 291 -543 483 -537
<< properties >>
string FIXED_BBOX -650 -658 650 658
string gencell sky130_fd_pr__nfet_g5v0d10v5
string library sky130
string parameters w 4.65 l 1.0 m 1 nf 4 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
