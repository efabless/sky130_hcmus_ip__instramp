magic
tech sky130A
magscale 1 2
timestamp 1717127936
<< dnwell >>
rect -60 -20 15946 3505
<< pwell >>
rect 15152 8984 20089 16096
rect 17204 -153 20102 85
rect 9975 -10266 10165 -329
<< locali >>
rect -285 16347 41 16348
rect -285 16021 20143 16347
rect -285 15400 41 16021
rect 154 15496 15034 15928
rect 15145 15400 20143 16021
rect -285 15200 20143 15400
rect -285 15000 41 15200
rect 15145 15192 20143 15200
rect 15145 15000 16535 15192
rect -285 14800 16535 15000
rect -285 14600 41 14800
rect 15145 14600 16535 14800
rect -285 14400 16535 14600
rect -285 14200 41 14400
rect 15145 14200 16535 14400
rect -285 14000 16535 14200
rect -285 13800 41 14000
rect 15145 13800 16535 14000
rect -285 13600 16535 13800
rect -285 13400 41 13600
rect 15145 13400 16535 13600
rect -285 13200 16535 13400
rect -285 12592 41 13200
rect 153 12652 15033 13084
rect 15145 12592 16535 13200
rect -285 12486 16535 12592
rect -285 11900 41 12486
rect 154 11994 15034 12426
rect 15145 11900 16535 12486
rect -285 11700 16535 11900
rect -285 11500 41 11700
rect 15145 11500 16535 11700
rect -285 11300 16535 11500
rect -285 11100 41 11300
rect 15145 11100 16535 11300
rect -285 10900 16535 11100
rect -285 10700 41 10900
rect 15145 10700 16535 10900
rect -285 10500 16535 10700
rect -285 10300 41 10500
rect 15145 10300 16535 10500
rect -285 10100 16535 10300
rect -285 9900 41 10100
rect 15145 9900 16535 10100
rect -285 9700 16535 9900
rect -285 9116 41 9700
rect 154 9150 15034 9582
rect 15145 9116 16535 9700
rect -285 9020 16535 9116
rect -285 -9044 -151 9020
rect -90 8722 90 8855
rect -90 4616 106 8722
rect 400 8000 1200 8800
rect 3077 5215 3274 8854
rect 3077 5125 3182 5215
rect 3272 5125 3274 5215
rect 3077 4617 3274 5125
rect 6260 4617 6457 8854
rect 9444 4617 9641 8854
rect 12629 4617 12826 8854
rect -90 -3815 43 4616
rect 77 4306 15816 4389
rect 77 4196 1313 4306
rect 3046 149 3317 4306
rect 6230 149 6501 4306
rect 9414 149 9685 4306
rect 12598 149 12869 4306
rect 77 54 15816 149
rect 16172 86 16534 9020
rect 16647 204 17080 15084
rect 17200 86 17400 15192
rect 17600 86 17800 15192
rect 18000 86 18200 15192
rect 18400 86 18600 15192
rect 18800 86 19000 15192
rect 19200 86 19400 15192
rect 19491 203 19924 15083
rect 20029 86 20143 15192
rect 16172 -130 20143 86
rect 195 -187 20143 -130
rect -90 -3915 -73 -3815
rect 27 -3915 43 -3815
rect -90 -8884 43 -3915
rect -90 -8984 -74 -8884
rect 26 -8984 43 -8884
rect -90 -8998 43 -8984
rect 126 -5114 194 -3642
rect 9940 -3745 10292 -187
rect 15916 -188 20143 -187
rect 10007 -3815 10136 -3800
rect 10007 -3915 10022 -3815
rect 10122 -3915 10136 -3815
rect 126 -5115 9956 -5114
rect 126 -5205 9845 -5115
rect 9935 -5205 9956 -5115
rect 126 -5211 9956 -5205
rect 126 -9044 194 -5211
rect 10007 -8883 10136 -3915
rect 10963 -5021 11093 -4830
rect 20029 -5092 20143 -188
rect 10223 -5115 20143 -5092
rect 10223 -5205 10246 -5115
rect 10336 -5205 20143 -5115
rect 10223 -5232 20143 -5205
rect 10007 -8983 10022 -8883
rect 10122 -8983 10136 -8883
rect 10007 -8998 10136 -8983
rect -285 -10160 194 -9044
rect 9933 -10160 10238 -9040
rect 20029 -10160 20143 -5232
rect -285 -10194 20143 -10160
rect -284 -10274 20143 -10194
<< viali >>
rect -73 -3915 27 -3815
rect -74 -8984 26 -8884
rect 10022 -3915 10122 -3815
rect 9845 -5205 9935 -5115
rect 10246 -5205 10336 -5115
rect 10236 -5743 10322 -5355
rect 10022 -8983 10122 -8883
<< metal1 >>
rect 154 15917 15034 15928
rect 154 15505 12735 15917
rect 12836 15505 15034 15917
rect 154 15496 15034 15505
rect 153 13073 15033 13084
rect 153 12660 9439 13073
rect 9681 12660 15033 13073
rect 153 12652 15033 12660
rect 154 11994 15034 12426
rect 4849 9765 4969 11994
rect 4849 9675 4865 9765
rect 4955 9675 4969 9765
rect 4849 9660 4969 9675
rect 154 9150 15034 9582
rect -461 5220 110 5230
rect -461 5120 0 5220
rect 100 5120 110 5220
rect -461 5110 110 5120
rect 1666 5015 1786 9150
rect 4849 9075 4969 9090
rect 4849 8985 4865 9075
rect 4955 8985 4969 9075
rect 1666 4935 1686 5015
rect 1766 4935 1786 5015
rect 1666 4924 1786 4935
rect 3166 5215 3286 5230
rect 3166 5125 3182 5215
rect 3272 5125 3286 5215
rect -461 4495 102 4615
rect 3166 4495 3286 5125
rect 4849 5080 4969 8985
rect 4849 5000 4870 5080
rect 4950 5000 4969 5080
rect 4849 4990 4969 5000
rect 12726 9078 12846 9090
rect 12726 8978 12736 9078
rect 12836 8978 12846 9078
rect 12726 4801 12846 8978
rect 16647 8844 17080 15084
rect 16647 8610 16660 8844
rect 17070 8610 17080 8844
rect 12726 4701 12735 4801
rect 12835 4701 12846 4801
rect 12726 4690 12846 4701
rect 13550 5280 13670 5290
rect 13550 5180 13560 5280
rect 13660 5180 13670 5280
rect 13550 4495 13670 5180
rect -10 812 110 4381
rect -256 692 110 812
rect -461 -618 -300 -607
rect -461 -678 -370 -618
rect -310 -678 -300 -618
rect -461 -687 -300 -678
rect -256 -4622 -136 692
rect 2909 446 3064 4125
rect 1530 405 1680 409
rect 1530 395 1564 405
rect 1530 297 1564 302
rect 1587 297 1680 405
rect 2909 377 3133 446
rect 2893 325 2980 377
rect 3117 325 3133 377
rect 1530 -405 1680 297
rect 3009 -295 3133 325
rect 3176 -33 3296 4384
rect 12726 4370 12846 4381
rect 12726 4270 12737 4370
rect 12837 4270 12846 4370
rect 6090 378 6245 4125
rect 6090 325 6158 378
rect 6230 325 6245 378
rect 3176 -123 3191 -33
rect 3281 -123 3296 -33
rect 3176 -139 3296 -123
rect 3009 -364 3061 -295
rect 7211 -424 7331 4234
rect 10393 151 10513 4234
rect 10393 20 10404 151
rect 10503 20 10513 151
rect 10393 10 10513 20
rect 12726 -35 12846 4270
rect 12726 -125 12741 -35
rect 12821 -125 12846 -35
rect 12726 -140 12846 -125
rect 13995 374 14416 409
rect 13995 322 14013 374
rect 14293 322 14416 374
rect 15639 377 15851 4125
rect 15639 325 15730 377
rect 15840 325 15851 377
rect 13995 -314 14416 322
rect 16647 204 17080 8610
rect 19491 5280 19924 15083
rect 19491 5180 19500 5280
rect 19914 5180 19924 5280
rect 19491 360 19924 5180
rect 20059 4030 20575 4043
rect 20059 3800 20070 4030
rect 20300 3800 20575 4030
rect 20059 3786 20575 3800
rect 19491 334 19925 360
rect 19491 214 20214 334
rect 5970 -3603 6123 -3580
rect 3523 -3642 3645 -3617
rect 3523 -3722 3546 -3642
rect 3626 -3722 3645 -3642
rect -90 -4038 140 -3958
rect -90 -4146 140 -4066
rect -90 -4254 140 -4174
rect -90 -4362 140 -4282
rect -90 -4470 140 -4390
rect -256 -4702 -10 -4622
rect 3523 -5132 3645 -3722
rect 5970 -3723 5987 -3603
rect 6107 -3723 6123 -3603
rect 3523 -5212 3547 -5132
rect 3627 -5212 3645 -5132
rect 3523 -5229 3645 -5212
rect 5970 -5563 6123 -3723
rect 12220 -3610 12340 -3600
rect 12220 -3710 12230 -3610
rect 12330 -3710 12340 -3610
rect 12220 -4613 12340 -3710
rect 12220 -4713 12230 -4613
rect 12330 -4713 12340 -4613
rect 12220 -4720 12340 -4713
rect 9830 -5115 9950 -5100
rect 9830 -5205 9845 -5115
rect 9935 -5205 9950 -5115
rect 9830 -5220 9950 -5205
rect 10223 -5115 10363 -5092
rect 10223 -5205 10246 -5115
rect 10336 -5205 10363 -5115
rect 10223 -5232 10363 -5205
rect 10223 -5355 10569 -5334
rect -461 -5755 -10 -5675
rect 10223 -5743 10236 -5355
rect 10322 -5743 10569 -5355
rect 10223 -5756 10569 -5743
rect -90 -6506 11093 -6500
rect -90 -6573 10970 -6506
rect 11087 -6573 11093 -6506
rect -90 -6580 11093 -6573
rect -90 -6646 11735 -6640
rect -90 -6713 11612 -6646
rect 11729 -6713 11735 -6646
rect -90 -6720 11735 -6713
rect -90 -6787 12627 -6780
rect -90 -6854 12504 -6787
rect 12621 -6854 12627 -6787
rect -90 -6860 12627 -6854
rect -90 -6926 14043 -6920
rect -90 -6993 13920 -6926
rect 14037 -6993 14043 -6926
rect -90 -7000 14043 -6993
rect -90 -7067 16486 -7060
rect -90 -7134 16363 -7067
rect 16480 -7134 16486 -7067
rect -90 -7140 16486 -7134
rect 866 -8705 996 -8690
rect 866 -8805 880 -8705
rect 980 -8805 996 -8705
rect -90 -9106 -10 -9026
rect 866 -9106 996 -8805
rect 1508 -8705 1638 -8690
rect 1508 -8805 1521 -8705
rect 1621 -8805 1638 -8705
rect 1508 -9030 1638 -8805
rect 2400 -8705 2530 -8690
rect 2400 -8805 2415 -8705
rect 2515 -8805 2530 -8705
rect 2400 -9060 2530 -8805
rect 3523 -8717 3646 -8707
rect 3523 -8817 3536 -8717
rect 3636 -8817 3646 -8717
rect -90 -9214 -10 -9134
rect -90 -9322 -10 -9242
rect -90 -9430 -10 -9350
rect -90 -9538 -10 -9458
rect 3523 -9697 3646 -8817
rect 3816 -8719 3946 -8707
rect 3816 -8819 3832 -8719
rect 3932 -8819 3946 -8719
rect 3816 -9007 3946 -8819
rect 6259 -8719 6389 -8710
rect 6259 -8819 6275 -8719
rect 6375 -8819 6389 -8719
rect 6259 -9006 6389 -8819
rect 3523 -9767 3550 -9697
rect 3620 -9767 3646 -9697
rect 20094 -9700 20214 214
rect 20094 -9760 20101 -9700
rect 20207 -9760 20214 -9700
rect 20094 -9766 20214 -9760
rect 3523 -9787 3646 -9767
<< via1 >>
rect 12735 15505 12836 15917
rect 9439 12660 9681 13073
rect 4865 9675 4955 9765
rect 0 5120 100 5220
rect 4865 8985 4955 9075
rect 1686 4935 1766 5015
rect 3182 5125 3272 5215
rect 4870 5000 4950 5080
rect 12736 8978 12836 9078
rect 16660 8610 17070 8844
rect 12735 4701 12835 4801
rect 13560 5180 13660 5280
rect 335 4275 425 4365
rect -370 -678 -310 -618
rect 1274 302 1564 395
rect 2980 325 3117 377
rect 3517 4276 3607 4366
rect 6700 4270 6790 4360
rect 9880 4270 9970 4360
rect 12737 4270 12837 4370
rect 4463 322 4755 374
rect 6158 325 6230 378
rect 3191 -123 3281 -33
rect 10404 20 10503 151
rect 12741 -125 12821 -35
rect 14013 322 14293 374
rect 15730 325 15840 377
rect 19500 5180 19914 5280
rect 20070 3800 20300 4030
rect -80 -676 -20 -616
rect 3546 -3722 3626 -3642
rect -73 -3915 27 -3815
rect 880 -4945 980 -4845
rect 1524 -4944 1624 -4844
rect 2415 -4946 2515 -4846
rect 5987 -3723 6107 -3603
rect 3830 -4945 3930 -4845
rect 3547 -5212 3627 -5132
rect 12230 -3710 12330 -3610
rect 10022 -3915 10122 -3815
rect 12230 -4713 12330 -4613
rect 6273 -4946 6373 -4846
rect 10979 -4945 11079 -4845
rect 11621 -4946 11721 -4846
rect 12513 -4946 12613 -4846
rect 13928 -4946 14028 -4846
rect 16370 -4946 16470 -4846
rect 9845 -5205 9935 -5115
rect 10246 -5205 10336 -5115
rect 10970 -6573 11087 -6506
rect 11612 -6713 11729 -6646
rect 12504 -6854 12621 -6787
rect 13920 -6993 14037 -6926
rect 16363 -7134 16480 -7067
rect 880 -8805 980 -8705
rect -74 -8984 26 -8884
rect 1521 -8805 1621 -8705
rect 2415 -8805 2515 -8705
rect 3536 -8817 3636 -8717
rect 3832 -8819 3932 -8719
rect 6275 -8819 6375 -8719
rect 10022 -8983 10122 -8883
rect 3550 -9767 3620 -9697
rect 20101 -9760 20207 -9700
<< metal2 >>
rect 12726 15917 12846 15928
rect 12726 15505 12735 15917
rect 12836 15505 12846 15917
rect 9431 13073 9691 13084
rect 9431 12660 9439 13073
rect 9681 12660 9691 13073
rect 4849 9765 4969 9780
rect 4849 9675 4865 9765
rect 4955 9675 4969 9765
rect 4849 9075 4969 9675
rect 4849 8985 4865 9075
rect 4955 8985 4969 9075
rect 4849 8970 4969 8985
rect 9431 8148 9691 12660
rect 12726 9078 12846 15505
rect 12726 8978 12736 9078
rect 12836 8978 12846 9078
rect 12726 8970 12846 8978
rect 12610 8844 17080 8857
rect 12610 8610 16660 8844
rect 17070 8610 17080 8844
rect 12610 8597 17080 8610
rect 12610 8148 12870 8597
rect 8772 7888 9691 8148
rect 11956 7888 12870 8148
rect 13550 5280 19924 5290
rect -10 5220 110 5230
rect -10 5120 0 5220
rect 100 5120 110 5220
rect -10 5110 110 5120
rect 600 5220 3286 5230
rect 600 5120 610 5220
rect 710 5215 3286 5220
rect 710 5125 3182 5215
rect 3272 5125 3286 5215
rect 13550 5180 13560 5280
rect 13660 5180 19500 5280
rect 19914 5180 19924 5280
rect 13550 5170 19924 5180
rect 710 5120 3286 5125
rect 600 5110 3286 5120
rect 4858 5080 4960 5090
rect 1675 5015 1779 5030
rect 1675 4935 1686 5015
rect 1766 4935 1779 5015
rect 1675 4372 1779 4935
rect 4858 5000 4870 5080
rect 4950 5000 4960 5080
rect 4858 4372 4960 5000
rect 327 4365 1779 4372
rect 327 4275 335 4365
rect 425 4275 1779 4365
rect 327 4268 1779 4275
rect 3510 4366 4960 4372
rect 12726 4801 12846 4810
rect 12726 4701 12735 4801
rect 12835 4701 12846 4801
rect 12726 4370 12846 4701
rect 3510 4276 3517 4366
rect 3607 4276 4960 4366
rect 3510 4270 4960 4276
rect 6690 4360 8983 4370
rect 6690 4270 6700 4360
rect 6790 4270 8983 4360
rect 6690 4260 8983 4270
rect 9871 4360 12149 4370
rect 9871 4270 9880 4360
rect 9970 4270 12149 4360
rect 9871 4261 12149 4270
rect 12726 4270 12737 4370
rect 12837 4270 12846 4370
rect 12726 4261 12846 4270
rect 15386 4030 20316 4043
rect 15386 3800 20070 4030
rect 20300 3800 20316 4030
rect 15386 3786 20316 3800
rect 1259 395 1680 409
rect 1259 302 1274 395
rect 1564 302 1680 395
rect 1259 291 1680 302
rect 1564 285 1680 291
rect 2903 377 3133 387
rect 2903 325 2980 377
rect 3117 325 3133 377
rect 2903 285 3133 325
rect 1564 169 3133 285
rect 4444 374 4864 410
rect 4444 322 4463 374
rect 4755 322 4864 374
rect 4444 284 4864 322
rect 6085 378 6239 396
rect 6085 325 6158 378
rect 6230 325 6239 378
rect 6085 284 6239 325
rect 13995 374 14416 409
rect 13995 322 14013 374
rect 14293 322 14416 374
rect 13995 284 14416 322
rect 15639 377 15850 387
rect 15639 325 15730 377
rect 15840 325 15850 377
rect 15639 284 15850 325
rect 4444 232 6304 284
rect 4707 163 6304 232
rect 13995 231 15850 284
rect 4707 151 10513 163
rect 4707 106 10404 151
rect 5970 20 10404 106
rect 10503 20 10513 151
rect 14219 106 15850 231
rect 5970 10 10513 20
rect 3176 -33 3645 -17
rect 3176 -123 3191 -33
rect 3281 -123 3645 -33
rect 3176 -139 3645 -123
rect -380 -616 -10 -607
rect -380 -618 -80 -616
rect -380 -678 -370 -618
rect -310 -676 -80 -618
rect -20 -676 -10 -616
rect -310 -678 -10 -676
rect -380 -687 -10 -678
rect 3523 -3642 3645 -139
rect 3523 -3722 3546 -3642
rect 3626 -3722 3645 -3642
rect 3523 -3733 3645 -3722
rect 5970 -3603 6123 10
rect 5970 -3723 5987 -3603
rect 6107 -3723 6123 -3603
rect 12220 -35 12836 -20
rect 12220 -125 12741 -35
rect 12821 -125 12836 -35
rect 12220 -140 12836 -125
rect 12220 -3610 12340 -140
rect 12220 -3710 12230 -3610
rect 12330 -3710 12340 -3610
rect 12220 -3720 12340 -3710
rect 5970 -3740 6123 -3723
rect -90 -3815 10136 -3800
rect -90 -3915 -73 -3815
rect 27 -3915 10022 -3815
rect 10122 -3915 10136 -3815
rect -90 -3930 10136 -3915
rect 12220 -4613 12340 -4606
rect 12220 -4713 12230 -4613
rect 12330 -4713 12340 -4613
rect 12220 -4720 12340 -4713
rect 866 -4845 996 -4830
rect 866 -4945 880 -4845
rect 980 -4945 996 -4845
rect 866 -8705 996 -4945
rect 866 -8805 880 -8705
rect 980 -8805 996 -8705
rect 866 -8820 996 -8805
rect 1508 -4844 1638 -4830
rect 1508 -4944 1524 -4844
rect 1624 -4944 1638 -4844
rect 1508 -8705 1638 -4944
rect 1508 -8805 1521 -8705
rect 1621 -8805 1638 -8705
rect 1508 -8820 1638 -8805
rect 2400 -4846 2530 -4830
rect 2400 -4946 2415 -4846
rect 2515 -4946 2530 -4846
rect 2400 -8705 2530 -4946
rect 3816 -4845 3946 -4830
rect 3816 -4945 3830 -4845
rect 3930 -4945 3946 -4845
rect 2400 -8805 2415 -8705
rect 2515 -8805 2530 -8705
rect 2400 -8820 2530 -8805
rect 3523 -5132 3646 -5117
rect 3523 -5212 3547 -5132
rect 3627 -5212 3646 -5132
rect 3523 -8717 3646 -5212
rect 3523 -8817 3536 -8717
rect 3636 -8817 3646 -8717
rect 3523 -8829 3646 -8817
rect 3816 -8719 3946 -4945
rect 3816 -8819 3832 -8719
rect 3932 -8819 3946 -8719
rect 3816 -8829 3946 -8819
rect 6259 -4846 6389 -4830
rect 6259 -4946 6273 -4846
rect 6373 -4946 6389 -4846
rect 6259 -8719 6389 -4946
rect 10963 -4845 11093 -4830
rect 10963 -4945 10979 -4845
rect 11079 -4945 11093 -4845
rect 9820 -5115 10363 -5092
rect 9820 -5205 9845 -5115
rect 9935 -5205 10246 -5115
rect 10336 -5205 10363 -5115
rect 9820 -5232 10363 -5205
rect 6259 -8819 6275 -8719
rect 6375 -8819 6389 -8719
rect 6259 -8829 6389 -8819
rect 10963 -6506 11093 -4945
rect 10963 -6573 10970 -6506
rect 11087 -6573 11093 -6506
rect -90 -8883 10136 -8868
rect -90 -8884 10022 -8883
rect -90 -8984 -74 -8884
rect 26 -8983 10022 -8884
rect 10122 -8983 10136 -8883
rect 26 -8984 10136 -8983
rect -90 -8998 10136 -8984
rect 10963 -9106 11093 -6573
rect 11605 -4846 11735 -4830
rect 11605 -4946 11621 -4846
rect 11721 -4946 11735 -4846
rect 11605 -6646 11735 -4946
rect 11605 -6713 11612 -6646
rect 11729 -6713 11735 -6646
rect 11605 -9214 11735 -6713
rect 12497 -4846 12627 -4830
rect 12497 -4946 12513 -4846
rect 12613 -4946 12627 -4846
rect 12497 -6787 12627 -4946
rect 12497 -6854 12504 -6787
rect 12621 -6854 12627 -6787
rect 12497 -9322 12627 -6854
rect 13913 -4846 14043 -4830
rect 13913 -4946 13928 -4846
rect 14028 -4946 14043 -4846
rect 13913 -6926 14043 -4946
rect 13913 -6993 13920 -6926
rect 14037 -6993 14043 -6926
rect 13913 -9430 14043 -6993
rect 16356 -4846 16486 -4830
rect 16356 -4946 16370 -4846
rect 16470 -4946 16486 -4846
rect 16356 -7067 16486 -4946
rect 16356 -7134 16363 -7067
rect 16480 -7134 16486 -7067
rect 16356 -9538 16486 -7134
rect 3541 -9697 3631 -9684
rect 3541 -9767 3550 -9697
rect 3620 -9767 3631 -9697
rect 19612 -9700 20214 -9694
rect 19612 -9760 20101 -9700
rect 20207 -9760 20214 -9700
rect 19612 -9766 20214 -9760
rect 3541 -9774 3631 -9767
<< via2 >>
rect 0 5120 100 5220
rect 610 5120 710 5220
<< metal3 >>
rect -10 5220 720 5230
rect -10 5120 0 5220
rect 100 5120 610 5220
rect 710 5120 720 5220
rect -10 5110 720 5120
use RB_array_20  x1
timestamp 1717127688
transform 1 0 -1780 0 1 -5002
box 1690 -194 11784 4950
use RB_array_20  x2
timestamp 1717127688
transform 1 0 -1780 0 1 -10070
box 1690 -194 11784 4950
use RB_array_20  x3
timestamp 1717127688
transform 1 0 8317 0 1 -5002
box 1690 -194 11784 4950
use opamp  x4
timestamp 1717127688
transform 1 0 -3828 0 1 -243
box 3810 247 7000 9177
use opamp  x5
timestamp 1717127688
transform 1 0 -644 0 1 -243
box 3810 247 7000 9177
use opamp  x6
timestamp 1717127688
transform 1 0 8908 0 1 -243
box 3810 247 7000 9177
use RB_array_20  x7
timestamp 1717127688
transform 1 0 8317 0 1 -10070
box 1690 -194 11784 4950
use opamp  x8
timestamp 1717127688
transform 1 0 2540 0 1 -243
box 3810 247 7000 9177
use opamp  x9
timestamp 1717127688
transform 1 0 5724 0 1 -243
box 3810 247 7000 9177
use sky130_fd_pr__res_high_po_0p69_WX3C5M  XR1
timestamp 1717127688
transform 1 0 7594 0 1 10788
box -7606 -1804 7606 1804
use sky130_fd_pr__res_high_po_0p69_WX3C5M  XR2
timestamp 1717127688
transform 0 1 18285 -1 0 7644
box -7606 -1804 7606 1804
use sky130_fd_pr__res_high_po_0p69_WX3C5M  XR4
timestamp 1717127688
transform 1 0 7594 0 1 14290
box -7606 -1804 7606 1804
<< labels >>
flabel space -12 12486 15200 16094 0 FreeSans 8000 0 0 0 XR4
flabel space -12 8984 15200 12592 0 FreeSans 8000 0 0 0 XR1
flabel space 16493 37 20101 15249 0 FreeSans 8000 0 0 0 XR2
flabel space -90 -10264 10004 -5120 0 FreeSans 8000 0 0 0 x2
flabel space 10007 -10265 20101 -5121 0 FreeSans 8000 0 0 0 x7
flabel space 10007 -5197 20101 -53 0 FreeSans 8000 0 0 0 x3
flabel space -90 -5196 10004 -52 0 FreeSans 8000 0 0 0 x1
flabel space 12718 4 15908 8934 0 FreeSans 8000 0 0 0 x6
flabel space 9534 4 12724 8934 0 FreeSans 8000 0 0 0 x9
flabel space 6350 4 9540 8934 0 FreeSans 8000 0 0 0 x8
flabel space 3166 4 6356 8934 0 FreeSans 8000 0 0 0 x5
flabel space -18 4 3172 8934 0 FreeSans 8000 0 0 0 x4
flabel locali 634 8272 1004 8630 0 FreeSans 4800 0 0 0 VDD
port 1 nsew
flabel metal1 -461 5110 -341 5230 0 FreeSans 4800 0 0 0 V1
port 4 nsew
flabel metal1 -461 4495 -341 4615 0 FreeSans 4800 0 0 0 V2
port 5 nsew
flabel metal1 -90 -4038 -10 -3958 0 FreeSans 960 0 0 0 D0
port 6 nsew
flabel metal1 -90 -4146 -10 -4066 0 FreeSans 960 0 0 0 D1
port 7 nsew
flabel metal1 -90 -4254 -10 -4174 0 FreeSans 960 0 0 0 D2
port 8 nsew
flabel metal1 -90 -4362 -10 -4282 0 FreeSans 960 0 0 0 D3
port 9 nsew
flabel metal1 -90 -4470 -10 -4390 0 FreeSans 960 0 0 0 D4
port 10 nsew
flabel metal1 -90 -6580 -10 -6500 0 FreeSans 960 0 0 0 D5
port 11 nsew
flabel metal1 -90 -6720 -10 -6640 0 FreeSans 960 0 0 0 D6
port 12 nsew
flabel metal1 -90 -6860 -10 -6780 0 FreeSans 960 0 0 0 D7
port 13 nsew
flabel metal1 -90 -7000 -10 -6920 0 FreeSans 960 0 0 0 D8
port 14 nsew
flabel metal1 -90 -7140 -10 -7060 0 FreeSans 960 0 0 0 D9
port 15 nsew
flabel metal1 -461 -687 -381 -607 0 FreeSans 4800 0 0 0 AVOUT1
port 16 nsew
flabel metal1 -461 -5755 -381 -5675 0 FreeSans 4800 0 0 0 AVOUT2
port 17 nsew
flabel metal1 20316 3786 20575 4043 0 FreeSans 4800 0 0 0 VOUT
port 18 nsew
flabel locali -250 -10240 -50 -10040 0 FreeSans 4800 0 0 0 G
port 3 nsew
flabel locali 86 57 166 137 0 FreeSans 4800 0 0 0 VSS
port 2 nsew
<< end >>
