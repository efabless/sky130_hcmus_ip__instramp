magic
tech sky130A
magscale 1 2
timestamp 1716878682
<< mvnmos >>
rect -100 8093 100 8893
rect -100 7199 100 7999
rect -100 6305 100 7105
rect -100 5411 100 6211
rect -100 4517 100 5317
rect -100 3623 100 4423
rect -100 2729 100 3529
rect -100 1835 100 2635
rect -100 941 100 1741
rect -100 47 100 847
rect -100 -847 100 -47
rect -100 -1741 100 -941
rect -100 -2635 100 -1835
rect -100 -3529 100 -2729
rect -100 -4423 100 -3623
rect -100 -5317 100 -4517
rect -100 -6211 100 -5411
rect -100 -7105 100 -6305
rect -100 -7999 100 -7199
rect -100 -8893 100 -8093
<< mvndiff >>
rect -158 8881 -100 8893
rect -158 8105 -146 8881
rect -112 8105 -100 8881
rect -158 8093 -100 8105
rect 100 8881 158 8893
rect 100 8105 112 8881
rect 146 8105 158 8881
rect 100 8093 158 8105
rect -158 7987 -100 7999
rect -158 7211 -146 7987
rect -112 7211 -100 7987
rect -158 7199 -100 7211
rect 100 7987 158 7999
rect 100 7211 112 7987
rect 146 7211 158 7987
rect 100 7199 158 7211
rect -158 7093 -100 7105
rect -158 6317 -146 7093
rect -112 6317 -100 7093
rect -158 6305 -100 6317
rect 100 7093 158 7105
rect 100 6317 112 7093
rect 146 6317 158 7093
rect 100 6305 158 6317
rect -158 6199 -100 6211
rect -158 5423 -146 6199
rect -112 5423 -100 6199
rect -158 5411 -100 5423
rect 100 6199 158 6211
rect 100 5423 112 6199
rect 146 5423 158 6199
rect 100 5411 158 5423
rect -158 5305 -100 5317
rect -158 4529 -146 5305
rect -112 4529 -100 5305
rect -158 4517 -100 4529
rect 100 5305 158 5317
rect 100 4529 112 5305
rect 146 4529 158 5305
rect 100 4517 158 4529
rect -158 4411 -100 4423
rect -158 3635 -146 4411
rect -112 3635 -100 4411
rect -158 3623 -100 3635
rect 100 4411 158 4423
rect 100 3635 112 4411
rect 146 3635 158 4411
rect 100 3623 158 3635
rect -158 3517 -100 3529
rect -158 2741 -146 3517
rect -112 2741 -100 3517
rect -158 2729 -100 2741
rect 100 3517 158 3529
rect 100 2741 112 3517
rect 146 2741 158 3517
rect 100 2729 158 2741
rect -158 2623 -100 2635
rect -158 1847 -146 2623
rect -112 1847 -100 2623
rect -158 1835 -100 1847
rect 100 2623 158 2635
rect 100 1847 112 2623
rect 146 1847 158 2623
rect 100 1835 158 1847
rect -158 1729 -100 1741
rect -158 953 -146 1729
rect -112 953 -100 1729
rect -158 941 -100 953
rect 100 1729 158 1741
rect 100 953 112 1729
rect 146 953 158 1729
rect 100 941 158 953
rect -158 835 -100 847
rect -158 59 -146 835
rect -112 59 -100 835
rect -158 47 -100 59
rect 100 835 158 847
rect 100 59 112 835
rect 146 59 158 835
rect 100 47 158 59
rect -158 -59 -100 -47
rect -158 -835 -146 -59
rect -112 -835 -100 -59
rect -158 -847 -100 -835
rect 100 -59 158 -47
rect 100 -835 112 -59
rect 146 -835 158 -59
rect 100 -847 158 -835
rect -158 -953 -100 -941
rect -158 -1729 -146 -953
rect -112 -1729 -100 -953
rect -158 -1741 -100 -1729
rect 100 -953 158 -941
rect 100 -1729 112 -953
rect 146 -1729 158 -953
rect 100 -1741 158 -1729
rect -158 -1847 -100 -1835
rect -158 -2623 -146 -1847
rect -112 -2623 -100 -1847
rect -158 -2635 -100 -2623
rect 100 -1847 158 -1835
rect 100 -2623 112 -1847
rect 146 -2623 158 -1847
rect 100 -2635 158 -2623
rect -158 -2741 -100 -2729
rect -158 -3517 -146 -2741
rect -112 -3517 -100 -2741
rect -158 -3529 -100 -3517
rect 100 -2741 158 -2729
rect 100 -3517 112 -2741
rect 146 -3517 158 -2741
rect 100 -3529 158 -3517
rect -158 -3635 -100 -3623
rect -158 -4411 -146 -3635
rect -112 -4411 -100 -3635
rect -158 -4423 -100 -4411
rect 100 -3635 158 -3623
rect 100 -4411 112 -3635
rect 146 -4411 158 -3635
rect 100 -4423 158 -4411
rect -158 -4529 -100 -4517
rect -158 -5305 -146 -4529
rect -112 -5305 -100 -4529
rect -158 -5317 -100 -5305
rect 100 -4529 158 -4517
rect 100 -5305 112 -4529
rect 146 -5305 158 -4529
rect 100 -5317 158 -5305
rect -158 -5423 -100 -5411
rect -158 -6199 -146 -5423
rect -112 -6199 -100 -5423
rect -158 -6211 -100 -6199
rect 100 -5423 158 -5411
rect 100 -6199 112 -5423
rect 146 -6199 158 -5423
rect 100 -6211 158 -6199
rect -158 -6317 -100 -6305
rect -158 -7093 -146 -6317
rect -112 -7093 -100 -6317
rect -158 -7105 -100 -7093
rect 100 -6317 158 -6305
rect 100 -7093 112 -6317
rect 146 -7093 158 -6317
rect 100 -7105 158 -7093
rect -158 -7211 -100 -7199
rect -158 -7987 -146 -7211
rect -112 -7987 -100 -7211
rect -158 -7999 -100 -7987
rect 100 -7211 158 -7199
rect 100 -7987 112 -7211
rect 146 -7987 158 -7211
rect 100 -7999 158 -7987
rect -158 -8105 -100 -8093
rect -158 -8881 -146 -8105
rect -112 -8881 -100 -8105
rect -158 -8893 -100 -8881
rect 100 -8105 158 -8093
rect 100 -8881 112 -8105
rect 146 -8881 158 -8105
rect 100 -8893 158 -8881
<< mvndiffc >>
rect -146 8105 -112 8881
rect 112 8105 146 8881
rect -146 7211 -112 7987
rect 112 7211 146 7987
rect -146 6317 -112 7093
rect 112 6317 146 7093
rect -146 5423 -112 6199
rect 112 5423 146 6199
rect -146 4529 -112 5305
rect 112 4529 146 5305
rect -146 3635 -112 4411
rect 112 3635 146 4411
rect -146 2741 -112 3517
rect 112 2741 146 3517
rect -146 1847 -112 2623
rect 112 1847 146 2623
rect -146 953 -112 1729
rect 112 953 146 1729
rect -146 59 -112 835
rect 112 59 146 835
rect -146 -835 -112 -59
rect 112 -835 146 -59
rect -146 -1729 -112 -953
rect 112 -1729 146 -953
rect -146 -2623 -112 -1847
rect 112 -2623 146 -1847
rect -146 -3517 -112 -2741
rect 112 -3517 146 -2741
rect -146 -4411 -112 -3635
rect 112 -4411 146 -3635
rect -146 -5305 -112 -4529
rect 112 -5305 146 -4529
rect -146 -6199 -112 -5423
rect 112 -6199 146 -5423
rect -146 -7093 -112 -6317
rect 112 -7093 146 -6317
rect -146 -7987 -112 -7211
rect 112 -7987 146 -7211
rect -146 -8881 -112 -8105
rect 112 -8881 146 -8105
<< poly >>
rect -100 8893 100 8919
rect -100 8067 100 8093
rect -100 7999 100 8025
rect -100 7173 100 7199
rect -100 7105 100 7131
rect -100 6279 100 6305
rect -100 6211 100 6237
rect -100 5385 100 5411
rect -100 5317 100 5343
rect -100 4491 100 4517
rect -100 4423 100 4449
rect -100 3597 100 3623
rect -100 3529 100 3555
rect -100 2703 100 2729
rect -100 2635 100 2661
rect -100 1809 100 1835
rect -100 1741 100 1767
rect -100 915 100 941
rect -100 847 100 873
rect -100 21 100 47
rect -100 -47 100 -21
rect -100 -873 100 -847
rect -100 -941 100 -915
rect -100 -1767 100 -1741
rect -100 -1835 100 -1809
rect -100 -2661 100 -2635
rect -100 -2729 100 -2703
rect -100 -3555 100 -3529
rect -100 -3623 100 -3597
rect -100 -4449 100 -4423
rect -100 -4517 100 -4491
rect -100 -5343 100 -5317
rect -100 -5411 100 -5385
rect -100 -6237 100 -6211
rect -100 -6305 100 -6279
rect -100 -7131 100 -7105
rect -100 -7199 100 -7173
rect -100 -8025 100 -7999
rect -100 -8093 100 -8067
rect -100 -8919 100 -8893
<< locali >>
rect -146 8881 -112 8897
rect -146 8089 -112 8105
rect 112 8881 146 8897
rect 112 8089 146 8105
rect -146 7987 -112 8003
rect -146 7195 -112 7211
rect 112 7987 146 8003
rect 112 7195 146 7211
rect -146 7093 -112 7109
rect -146 6301 -112 6317
rect 112 7093 146 7109
rect 112 6301 146 6317
rect -146 6199 -112 6215
rect -146 5407 -112 5423
rect 112 6199 146 6215
rect 112 5407 146 5423
rect -146 5305 -112 5321
rect -146 4513 -112 4529
rect 112 5305 146 5321
rect 112 4513 146 4529
rect -146 4411 -112 4427
rect -146 3619 -112 3635
rect 112 4411 146 4427
rect 112 3619 146 3635
rect -146 3517 -112 3533
rect -146 2725 -112 2741
rect 112 3517 146 3533
rect 112 2725 146 2741
rect -146 2623 -112 2639
rect -146 1831 -112 1847
rect 112 2623 146 2639
rect 112 1831 146 1847
rect -146 1729 -112 1745
rect -146 937 -112 953
rect 112 1729 146 1745
rect 112 937 146 953
rect -146 835 -112 851
rect -146 43 -112 59
rect 112 835 146 851
rect 112 43 146 59
rect -146 -59 -112 -43
rect -146 -851 -112 -835
rect 112 -59 146 -43
rect 112 -851 146 -835
rect -146 -953 -112 -937
rect -146 -1745 -112 -1729
rect 112 -953 146 -937
rect 112 -1745 146 -1729
rect -146 -1847 -112 -1831
rect -146 -2639 -112 -2623
rect 112 -1847 146 -1831
rect 112 -2639 146 -2623
rect -146 -2741 -112 -2725
rect -146 -3533 -112 -3517
rect 112 -2741 146 -2725
rect 112 -3533 146 -3517
rect -146 -3635 -112 -3619
rect -146 -4427 -112 -4411
rect 112 -3635 146 -3619
rect 112 -4427 146 -4411
rect -146 -4529 -112 -4513
rect -146 -5321 -112 -5305
rect 112 -4529 146 -4513
rect 112 -5321 146 -5305
rect -146 -5423 -112 -5407
rect -146 -6215 -112 -6199
rect 112 -5423 146 -5407
rect 112 -6215 146 -6199
rect -146 -6317 -112 -6301
rect -146 -7109 -112 -7093
rect 112 -6317 146 -6301
rect 112 -7109 146 -7093
rect -146 -7211 -112 -7195
rect -146 -8003 -112 -7987
rect 112 -7211 146 -7195
rect 112 -8003 146 -7987
rect -146 -8105 -112 -8089
rect -146 -8897 -112 -8881
rect 112 -8105 146 -8089
rect 112 -8897 146 -8881
<< viali >>
rect -146 8105 -112 8881
rect 112 8105 146 8881
rect -146 7211 -112 7987
rect 112 7211 146 7987
rect -146 6317 -112 7093
rect 112 6317 146 7093
rect -146 5423 -112 6199
rect 112 5423 146 6199
rect -146 4529 -112 5305
rect 112 4529 146 5305
rect -146 3635 -112 4411
rect 112 3635 146 4411
rect -146 2741 -112 3517
rect 112 2741 146 3517
rect -146 1847 -112 2623
rect 112 1847 146 2623
rect -146 953 -112 1729
rect 112 953 146 1729
rect -146 59 -112 835
rect 112 59 146 835
rect -146 -835 -112 -59
rect 112 -835 146 -59
rect -146 -1729 -112 -953
rect 112 -1729 146 -953
rect -146 -2623 -112 -1847
rect 112 -2623 146 -1847
rect -146 -3517 -112 -2741
rect 112 -3517 146 -2741
rect -146 -4411 -112 -3635
rect 112 -4411 146 -3635
rect -146 -5305 -112 -4529
rect 112 -5305 146 -4529
rect -146 -6199 -112 -5423
rect 112 -6199 146 -5423
rect -146 -7093 -112 -6317
rect 112 -7093 146 -6317
rect -146 -7987 -112 -7211
rect 112 -7987 146 -7211
rect -146 -8881 -112 -8105
rect 112 -8881 146 -8105
<< metal1 >>
rect -152 8881 -106 8893
rect -152 8105 -146 8881
rect -112 8105 -106 8881
rect -152 8093 -106 8105
rect 106 8881 152 8893
rect 106 8105 112 8881
rect 146 8105 152 8881
rect 106 8093 152 8105
rect -152 7987 -106 7999
rect -152 7211 -146 7987
rect -112 7211 -106 7987
rect -152 7199 -106 7211
rect 106 7987 152 7999
rect 106 7211 112 7987
rect 146 7211 152 7987
rect 106 7199 152 7211
rect -152 7093 -106 7105
rect -152 6317 -146 7093
rect -112 6317 -106 7093
rect -152 6305 -106 6317
rect 106 7093 152 7105
rect 106 6317 112 7093
rect 146 6317 152 7093
rect 106 6305 152 6317
rect -152 6199 -106 6211
rect -152 5423 -146 6199
rect -112 5423 -106 6199
rect -152 5411 -106 5423
rect 106 6199 152 6211
rect 106 5423 112 6199
rect 146 5423 152 6199
rect 106 5411 152 5423
rect -152 5305 -106 5317
rect -152 4529 -146 5305
rect -112 4529 -106 5305
rect -152 4517 -106 4529
rect 106 5305 152 5317
rect 106 4529 112 5305
rect 146 4529 152 5305
rect 106 4517 152 4529
rect -152 4411 -106 4423
rect -152 3635 -146 4411
rect -112 3635 -106 4411
rect -152 3623 -106 3635
rect 106 4411 152 4423
rect 106 3635 112 4411
rect 146 3635 152 4411
rect 106 3623 152 3635
rect -152 3517 -106 3529
rect -152 2741 -146 3517
rect -112 2741 -106 3517
rect -152 2729 -106 2741
rect 106 3517 152 3529
rect 106 2741 112 3517
rect 146 2741 152 3517
rect 106 2729 152 2741
rect -152 2623 -106 2635
rect -152 1847 -146 2623
rect -112 1847 -106 2623
rect -152 1835 -106 1847
rect 106 2623 152 2635
rect 106 1847 112 2623
rect 146 1847 152 2623
rect 106 1835 152 1847
rect -152 1729 -106 1741
rect -152 953 -146 1729
rect -112 953 -106 1729
rect -152 941 -106 953
rect 106 1729 152 1741
rect 106 953 112 1729
rect 146 953 152 1729
rect 106 941 152 953
rect -152 835 -106 847
rect -152 59 -146 835
rect -112 59 -106 835
rect -152 47 -106 59
rect 106 835 152 847
rect 106 59 112 835
rect 146 59 152 835
rect 106 47 152 59
rect -152 -59 -106 -47
rect -152 -835 -146 -59
rect -112 -835 -106 -59
rect -152 -847 -106 -835
rect 106 -59 152 -47
rect 106 -835 112 -59
rect 146 -835 152 -59
rect 106 -847 152 -835
rect -152 -953 -106 -941
rect -152 -1729 -146 -953
rect -112 -1729 -106 -953
rect -152 -1741 -106 -1729
rect 106 -953 152 -941
rect 106 -1729 112 -953
rect 146 -1729 152 -953
rect 106 -1741 152 -1729
rect -152 -1847 -106 -1835
rect -152 -2623 -146 -1847
rect -112 -2623 -106 -1847
rect -152 -2635 -106 -2623
rect 106 -1847 152 -1835
rect 106 -2623 112 -1847
rect 146 -2623 152 -1847
rect 106 -2635 152 -2623
rect -152 -2741 -106 -2729
rect -152 -3517 -146 -2741
rect -112 -3517 -106 -2741
rect -152 -3529 -106 -3517
rect 106 -2741 152 -2729
rect 106 -3517 112 -2741
rect 146 -3517 152 -2741
rect 106 -3529 152 -3517
rect -152 -3635 -106 -3623
rect -152 -4411 -146 -3635
rect -112 -4411 -106 -3635
rect -152 -4423 -106 -4411
rect 106 -3635 152 -3623
rect 106 -4411 112 -3635
rect 146 -4411 152 -3635
rect 106 -4423 152 -4411
rect -152 -4529 -106 -4517
rect -152 -5305 -146 -4529
rect -112 -5305 -106 -4529
rect -152 -5317 -106 -5305
rect 106 -4529 152 -4517
rect 106 -5305 112 -4529
rect 146 -5305 152 -4529
rect 106 -5317 152 -5305
rect -152 -5423 -106 -5411
rect -152 -6199 -146 -5423
rect -112 -6199 -106 -5423
rect -152 -6211 -106 -6199
rect 106 -5423 152 -5411
rect 106 -6199 112 -5423
rect 146 -6199 152 -5423
rect 106 -6211 152 -6199
rect -152 -6317 -106 -6305
rect -152 -7093 -146 -6317
rect -112 -7093 -106 -6317
rect -152 -7105 -106 -7093
rect 106 -6317 152 -6305
rect 106 -7093 112 -6317
rect 146 -7093 152 -6317
rect 106 -7105 152 -7093
rect -152 -7211 -106 -7199
rect -152 -7987 -146 -7211
rect -112 -7987 -106 -7211
rect -152 -7999 -106 -7987
rect 106 -7211 152 -7199
rect 106 -7987 112 -7211
rect 146 -7987 152 -7211
rect 106 -7999 152 -7987
rect -152 -8105 -106 -8093
rect -152 -8881 -146 -8105
rect -112 -8881 -106 -8105
rect -152 -8893 -106 -8881
rect 106 -8105 152 -8093
rect 106 -8881 112 -8105
rect 146 -8881 152 -8105
rect 106 -8893 152 -8881
<< properties >>
string gencell sky130_fd_pr__nfet_g5v0d10v5
string library sky130
string parameters w 4.0 l 1.0 m 20 nf 1 diffcov 100 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 0 botc 0 poverlap 0 doverlap 0 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 0 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
