* SPICE3 file created from IA_v4.ext - technology: sky130A

.subckt sky130_fd_pr__res_high_po_0p69_JKKHRG a_n199_n1768# a_n69_1206# a_n69_n1638#
X0 a_n69_1206# a_n69_n1638# a_n199_n1768# sky130_fd_pr__res_high_po_0p69 l=12.1
C0 a_n69_n1638# a_n199_n1768# 0.675f
C1 a_n69_1206# a_n199_n1768# 0.675f
.ends

.subckt sky130_fd_pr__res_high_po_0p69_Z3RMRJ a_48_1206# a_n186_n1638# a_n186_1206#
+ a_n316_n1768# a_48_n1638#
X0 a_48_1206# a_48_n1638# a_n316_n1768# sky130_fd_pr__res_high_po_0p69 l=12.1
X1 a_n186_1206# a_n186_n1638# a_n316_n1768# sky130_fd_pr__res_high_po_0p69 l=12.1
C0 a_n186_1206# a_48_1206# 0.296f
C1 a_n186_n1638# a_48_n1638# 0.296f
C2 a_48_n1638# a_n316_n1768# 0.465f
C3 a_48_1206# a_n316_n1768# 0.465f
C4 a_n186_n1638# a_n316_n1768# 0.465f
C5 a_n186_1206# a_n316_n1768# 0.465f
.ends

.subckt sky130_fd_pr__res_high_po_0p69_Z3RMR6 a_516_n1638# a_48_1206# a_n654_1206#
+ a_n888_1206# a_n186_n1638# a_n186_1206# a_750_1206# a_n654_n1638# a_282_1206# a_282_n1638#
+ a_48_n1638# a_750_n1638# a_n420_n1638# a_516_1206# a_n1018_n1768# a_n420_1206# a_n888_n1638#
X0 a_n420_1206# a_n420_n1638# a_n1018_n1768# sky130_fd_pr__res_high_po_0p69 l=12.1
X1 a_48_1206# a_48_n1638# a_n1018_n1768# sky130_fd_pr__res_high_po_0p69 l=12.1
X2 a_750_1206# a_750_n1638# a_n1018_n1768# sky130_fd_pr__res_high_po_0p69 l=12.1
X3 a_n888_1206# a_n888_n1638# a_n1018_n1768# sky130_fd_pr__res_high_po_0p69 l=12.1
X4 a_282_1206# a_282_n1638# a_n1018_n1768# sky130_fd_pr__res_high_po_0p69 l=12.1
X5 a_n654_1206# a_n654_n1638# a_n1018_n1768# sky130_fd_pr__res_high_po_0p69 l=12.1
X6 a_n186_1206# a_n186_n1638# a_n1018_n1768# sky130_fd_pr__res_high_po_0p69 l=12.1
X7 a_516_1206# a_516_n1638# a_n1018_n1768# sky130_fd_pr__res_high_po_0p69 l=12.1
C0 a_n420_n1638# a_n654_n1638# 0.296f
C1 a_48_n1638# a_n186_n1638# 0.296f
C2 a_n888_1206# a_n654_1206# 0.296f
C3 a_282_1206# a_516_1206# 0.296f
C4 a_n186_1206# a_48_1206# 0.296f
C5 a_48_n1638# a_282_n1638# 0.296f
C6 a_n420_1206# a_n654_1206# 0.296f
C7 a_750_1206# a_516_1206# 0.296f
C8 a_n888_n1638# a_n654_n1638# 0.296f
C9 a_n420_1206# a_n186_1206# 0.296f
C10 a_n420_n1638# a_n186_n1638# 0.296f
C11 a_516_n1638# a_750_n1638# 0.296f
C12 a_516_n1638# a_282_n1638# 0.296f
C13 a_282_1206# a_48_1206# 0.296f
C14 a_750_n1638# a_n1018_n1768# 0.465f
C15 a_750_1206# a_n1018_n1768# 0.465f
C16 a_516_n1638# a_n1018_n1768# 0.255f
C17 a_516_1206# a_n1018_n1768# 0.255f
C18 a_282_n1638# a_n1018_n1768# 0.255f
C19 a_282_1206# a_n1018_n1768# 0.255f
C20 a_48_n1638# a_n1018_n1768# 0.255f
C21 a_48_1206# a_n1018_n1768# 0.255f
C22 a_n186_n1638# a_n1018_n1768# 0.255f
C23 a_n186_1206# a_n1018_n1768# 0.255f
C24 a_n420_n1638# a_n1018_n1768# 0.255f
C25 a_n420_1206# a_n1018_n1768# 0.255f
C26 a_n654_n1638# a_n1018_n1768# 0.255f
C27 a_n654_1206# a_n1018_n1768# 0.255f
C28 a_n888_n1638# a_n1018_n1768# 0.465f
C29 a_n888_1206# a_n1018_n1768# 0.465f
.ends

.subckt sky130_fd_pr__res_high_po_0p69_YMHKRJ a_48_1206# a_n550_n1768# a_n186_n1638#
+ a_n186_1206# a_282_1206# a_282_n1638# a_48_n1638# a_n420_n1638# a_n420_1206#
X0 a_n420_1206# a_n420_n1638# a_n550_n1768# sky130_fd_pr__res_high_po_0p69 l=12.1
X1 a_48_1206# a_48_n1638# a_n550_n1768# sky130_fd_pr__res_high_po_0p69 l=12.1
X2 a_282_1206# a_282_n1638# a_n550_n1768# sky130_fd_pr__res_high_po_0p69 l=12.1
X3 a_n186_1206# a_n186_n1638# a_n550_n1768# sky130_fd_pr__res_high_po_0p69 l=12.1
C0 a_48_1206# a_282_1206# 0.296f
C1 a_48_n1638# a_282_n1638# 0.296f
C2 a_n186_1206# a_48_1206# 0.296f
C3 a_n186_1206# a_n420_1206# 0.296f
C4 a_n420_n1638# a_n186_n1638# 0.296f
C5 a_48_n1638# a_n186_n1638# 0.296f
C6 a_282_n1638# a_n550_n1768# 0.465f
C7 a_282_1206# a_n550_n1768# 0.465f
C8 a_48_n1638# a_n550_n1768# 0.255f
C9 a_48_1206# a_n550_n1768# 0.255f
C10 a_n186_n1638# a_n550_n1768# 0.255f
C11 a_n186_1206# a_n550_n1768# 0.255f
C12 a_n420_n1638# a_n550_n1768# 0.465f
C13 a_n420_1206# a_n550_n1768# 0.465f
.ends

.subckt sky130_fd_pr__res_high_po_0p69_HBQF5Z a_516_n1638# a_48_1206# a_n654_1206#
+ a_n888_1206# a_1452_1206# a_n1122_n1638# a_1452_n1638# a_n186_n1638# a_n186_1206#
+ a_n1954_n1768# a_1686_1206# a_750_1206# a_n654_n1638# a_n1590_1206# a_984_n1638#
+ a_984_1206# a_n1824_1206# a_n1590_n1638# a_1218_n1638# a_282_1206# a_n1122_1206#
+ a_1218_1206# a_282_n1638# a_48_n1638# a_750_n1638# a_n420_n1638# a_n1356_1206# a_516_1206#
+ a_n1356_n1638# a_1686_n1638# a_n420_1206# a_n1824_n1638# a_n888_n1638#
X0 a_n420_1206# a_n420_n1638# a_n1954_n1768# sky130_fd_pr__res_high_po_0p69 l=12.1
X1 a_1452_1206# a_1452_n1638# a_n1954_n1768# sky130_fd_pr__res_high_po_0p69 l=12.1
X2 a_n1824_1206# a_n1824_n1638# a_n1954_n1768# sky130_fd_pr__res_high_po_0p69 l=12.1
X3 a_n1590_1206# a_n1590_n1638# a_n1954_n1768# sky130_fd_pr__res_high_po_0p69 l=12.1
X4 a_48_1206# a_48_n1638# a_n1954_n1768# sky130_fd_pr__res_high_po_0p69 l=12.1
X5 a_984_1206# a_984_n1638# a_n1954_n1768# sky130_fd_pr__res_high_po_0p69 l=12.1
X6 a_n1356_1206# a_n1356_n1638# a_n1954_n1768# sky130_fd_pr__res_high_po_0p69 l=12.1
X7 a_1218_1206# a_1218_n1638# a_n1954_n1768# sky130_fd_pr__res_high_po_0p69 l=12.1
X8 a_750_1206# a_750_n1638# a_n1954_n1768# sky130_fd_pr__res_high_po_0p69 l=12.1
X9 a_n1122_1206# a_n1122_n1638# a_n1954_n1768# sky130_fd_pr__res_high_po_0p69 l=12.1
X10 a_n888_1206# a_n888_n1638# a_n1954_n1768# sky130_fd_pr__res_high_po_0p69 l=12.1
X11 a_282_1206# a_282_n1638# a_n1954_n1768# sky130_fd_pr__res_high_po_0p69 l=12.1
X12 a_n654_1206# a_n654_n1638# a_n1954_n1768# sky130_fd_pr__res_high_po_0p69 l=12.1
X13 a_n186_1206# a_n186_n1638# a_n1954_n1768# sky130_fd_pr__res_high_po_0p69 l=12.1
X14 a_516_1206# a_516_n1638# a_n1954_n1768# sky130_fd_pr__res_high_po_0p69 l=12.1
X15 a_1686_1206# a_1686_n1638# a_n1954_n1768# sky130_fd_pr__res_high_po_0p69 l=12.1
C0 a_1686_n1638# a_1452_n1638# 0.296f
C1 a_48_n1638# a_n186_n1638# 0.296f
C2 a_984_1206# a_1218_1206# 0.296f
C3 a_1452_1206# a_1218_1206# 0.296f
C4 a_750_1206# a_516_1206# 0.296f
C5 a_48_1206# a_282_1206# 0.296f
C6 a_n654_1206# a_n420_1206# 0.296f
C7 a_n1356_n1638# a_n1590_n1638# 0.296f
C8 a_n1122_n1638# a_n888_n1638# 0.296f
C9 a_n186_1206# a_n420_1206# 0.296f
C10 a_n1824_1206# a_n1590_1206# 0.296f
C11 a_n1824_n1638# a_n1590_n1638# 0.296f
C12 a_n888_n1638# a_n654_n1638# 0.296f
C13 a_1686_1206# a_1452_1206# 0.296f
C14 a_1452_n1638# a_1218_n1638# 0.296f
C15 a_516_1206# a_282_1206# 0.296f
C16 a_750_n1638# a_516_n1638# 0.296f
C17 a_48_1206# a_n186_1206# 0.296f
C18 a_n1356_1206# a_n1122_1206# 0.296f
C19 a_516_n1638# a_282_n1638# 0.296f
C20 a_n1356_n1638# a_n1122_n1638# 0.296f
C21 a_n420_n1638# a_n654_n1638# 0.296f
C22 a_n420_n1638# a_n186_n1638# 0.296f
C23 a_750_1206# a_984_1206# 0.296f
C24 a_48_n1638# a_282_n1638# 0.296f
C25 a_n888_1206# a_n654_1206# 0.296f
C26 a_n888_1206# a_n1122_1206# 0.296f
C27 a_984_n1638# a_1218_n1638# 0.296f
C28 a_n1590_1206# a_n1356_1206# 0.296f
C29 a_750_n1638# a_984_n1638# 0.296f
C30 a_1686_n1638# a_n1954_n1768# 0.465f
C31 a_1686_1206# a_n1954_n1768# 0.465f
C32 a_1452_n1638# a_n1954_n1768# 0.255f
C33 a_1452_1206# a_n1954_n1768# 0.255f
C34 a_1218_n1638# a_n1954_n1768# 0.255f
C35 a_1218_1206# a_n1954_n1768# 0.255f
C36 a_984_n1638# a_n1954_n1768# 0.255f
C37 a_984_1206# a_n1954_n1768# 0.255f
C38 a_750_n1638# a_n1954_n1768# 0.255f
C39 a_750_1206# a_n1954_n1768# 0.255f
C40 a_516_n1638# a_n1954_n1768# 0.255f
C41 a_516_1206# a_n1954_n1768# 0.255f
C42 a_282_n1638# a_n1954_n1768# 0.255f
C43 a_282_1206# a_n1954_n1768# 0.255f
C44 a_48_n1638# a_n1954_n1768# 0.255f
C45 a_48_1206# a_n1954_n1768# 0.255f
C46 a_n186_n1638# a_n1954_n1768# 0.255f
C47 a_n186_1206# a_n1954_n1768# 0.255f
C48 a_n420_n1638# a_n1954_n1768# 0.255f
C49 a_n420_1206# a_n1954_n1768# 0.255f
C50 a_n654_n1638# a_n1954_n1768# 0.255f
C51 a_n654_1206# a_n1954_n1768# 0.255f
C52 a_n888_n1638# a_n1954_n1768# 0.255f
C53 a_n888_1206# a_n1954_n1768# 0.255f
C54 a_n1122_n1638# a_n1954_n1768# 0.255f
C55 a_n1122_1206# a_n1954_n1768# 0.255f
C56 a_n1356_n1638# a_n1954_n1768# 0.255f
C57 a_n1356_1206# a_n1954_n1768# 0.255f
C58 a_n1590_n1638# a_n1954_n1768# 0.255f
C59 a_n1590_1206# a_n1954_n1768# 0.255f
C60 a_n1824_n1638# a_n1954_n1768# 0.465f
C61 a_n1824_1206# a_n1954_n1768# 0.465f
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_727CUP a_n100_n565# a_100_n477# a_n292_n699#
+ a_n158_n477#
X0 a_100_n477# a_n100_n565# a_n158_n477# a_n292_n699# sky130_fd_pr__nfet_g5v0d10v5 ad=1.38 pd=10.1 as=1.38 ps=10.1 w=4.77 l=1
C0 a_n158_n477# a_n100_n565# 0.107f
C1 a_100_n477# a_n100_n565# 0.107f
C2 a_100_n477# a_n158_n477# 0.261f
C3 a_100_n477# a_n292_n699# 0.53f
C4 a_n158_n477# a_n292_n699# 0.53f
C5 a_n100_n565# a_n292_n699# 0.714f
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_VU5C5A a_n287_n487# a_n421_n709# a_n229_n575#
+ a_229_n487# a_n29_n487# a_29_n575#
X0 a_229_n487# a_29_n575# a_n29_n487# a_n421_n709# sky130_fd_pr__nfet_g5v0d10v5 ad=1.41 pd=10.3 as=0.706 ps=5.16 w=4.87 l=1
X1 a_n29_n487# a_n229_n575# a_n287_n487# a_n421_n709# sky130_fd_pr__nfet_g5v0d10v5 ad=0.706 pd=5.16 as=1.41 ps=10.3 w=4.87 l=1
C0 a_29_n575# a_n229_n575# 0.104f
C1 a_n29_n487# a_29_n575# 0.11f
C2 a_n287_n487# a_n229_n575# 0.11f
C3 a_n287_n487# a_n29_n487# 0.267f
C4 a_229_n487# a_29_n575# 0.11f
C5 a_n29_n487# a_n229_n575# 0.11f
C6 a_229_n487# a_n29_n487# 0.267f
C7 a_229_n487# a_n421_n709# 0.54f
C8 a_n29_n487# a_n421_n709# 0.163f
C9 a_n287_n487# a_n421_n709# 0.54f
C10 a_29_n575# a_n421_n709# 0.651f
C11 a_n229_n575# a_n421_n709# 0.651f
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_J97EKB a_487_n438# a_n803_n438# a_29_n526# a_n745_n526#
+ a_n287_n438# a_n1061_n438# a_803_n526# a_745_n438# a_n229_n526# a_287_n526# a_n1003_n526#
+ a_229_n438# a_n545_n438# a_1003_n438# a_n487_n526# a_n1195_n660# a_545_n526# a_n29_n438#
X0 a_1003_n438# a_803_n526# a_745_n438# a_n1195_n660# sky130_fd_pr__nfet_g5v0d10v5 ad=1.27 pd=9.34 as=0.635 ps=4.67 w=4.38 l=1
X1 a_745_n438# a_545_n526# a_487_n438# a_n1195_n660# sky130_fd_pr__nfet_g5v0d10v5 ad=0.635 pd=4.67 as=0.635 ps=4.67 w=4.38 l=1
X2 a_487_n438# a_287_n526# a_229_n438# a_n1195_n660# sky130_fd_pr__nfet_g5v0d10v5 ad=0.635 pd=4.67 as=0.635 ps=4.67 w=4.38 l=1
X3 a_229_n438# a_29_n526# a_n29_n438# a_n1195_n660# sky130_fd_pr__nfet_g5v0d10v5 ad=0.635 pd=4.67 as=0.635 ps=4.67 w=4.38 l=1
X4 a_n29_n438# a_n229_n526# a_n287_n438# a_n1195_n660# sky130_fd_pr__nfet_g5v0d10v5 ad=0.635 pd=4.67 as=0.635 ps=4.67 w=4.38 l=1
X5 a_n545_n438# a_n745_n526# a_n803_n438# a_n1195_n660# sky130_fd_pr__nfet_g5v0d10v5 ad=0.635 pd=4.67 as=0.635 ps=4.67 w=4.38 l=1
X6 a_n287_n438# a_n487_n526# a_n545_n438# a_n1195_n660# sky130_fd_pr__nfet_g5v0d10v5 ad=0.635 pd=4.67 as=0.635 ps=4.67 w=4.38 l=1
X7 a_n803_n438# a_n1003_n526# a_n1061_n438# a_n1195_n660# sky130_fd_pr__nfet_g5v0d10v5 ad=0.635 pd=4.67 as=1.27 ps=9.34 w=4.38 l=1
C0 a_n745_n526# a_n1003_n526# 0.104f
C1 a_287_n526# a_487_n438# 0.099f
C2 a_1003_n438# a_803_n526# 0.099f
C3 a_n1061_n438# a_n803_n438# 0.24f
C4 a_29_n526# a_n29_n438# 0.099f
C5 a_487_n438# a_229_n438# 0.24f
C6 a_n487_n526# a_n545_n438# 0.099f
C7 a_745_n438# a_545_n526# 0.099f
C8 a_803_n526# a_745_n438# 0.099f
C9 a_n803_n438# a_n745_n526# 0.099f
C10 a_n545_n438# a_n287_n438# 0.24f
C11 a_n29_n438# a_229_n438# 0.24f
C12 a_n487_n526# a_n229_n526# 0.104f
C13 a_803_n526# a_545_n526# 0.104f
C14 a_n487_n526# a_n287_n438# 0.099f
C15 a_287_n526# a_29_n526# 0.104f
C16 a_n803_n438# a_n545_n438# 0.24f
C17 a_287_n526# a_545_n526# 0.104f
C18 a_29_n526# a_229_n438# 0.099f
C19 a_745_n438# a_487_n438# 0.24f
C20 a_n229_n526# a_n287_n438# 0.099f
C21 a_n1061_n438# a_n1003_n526# 0.099f
C22 a_n803_n438# a_n1003_n526# 0.099f
C23 a_1003_n438# a_745_n438# 0.24f
C24 a_n229_n526# a_n29_n438# 0.099f
C25 a_n29_n438# a_n287_n438# 0.24f
C26 a_487_n438# a_545_n526# 0.099f
C27 a_287_n526# a_229_n438# 0.099f
C28 a_n545_n438# a_n745_n526# 0.099f
C29 a_n487_n526# a_n745_n526# 0.104f
C30 a_29_n526# a_n229_n526# 0.104f
C31 a_1003_n438# a_n1195_n660# 0.489f
C32 a_745_n438# a_n1195_n660# 0.149f
C33 a_487_n438# a_n1195_n660# 0.149f
C34 a_229_n438# a_n1195_n660# 0.149f
C35 a_n29_n438# a_n1195_n660# 0.149f
C36 a_n287_n438# a_n1195_n660# 0.149f
C37 a_n545_n438# a_n1195_n660# 0.149f
C38 a_n803_n438# a_n1195_n660# 0.149f
C39 a_n1061_n438# a_n1195_n660# 0.489f
C40 a_803_n526# a_n1195_n660# 0.65f
C41 a_545_n526# a_n1195_n660# 0.587f
C42 a_287_n526# a_n1195_n660# 0.587f
C43 a_29_n526# a_n1195_n660# 0.587f
C44 a_n229_n526# a_n1195_n660# 0.587f
C45 a_n487_n526# a_n1195_n660# 0.587f
C46 a_n745_n526# a_n1195_n660# 0.587f
C47 a_n1003_n526# a_n1195_n660# 0.65f
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_S7E57E a_n229_n553# a_287_n553# a_229_n465# a_n545_n465#
+ a_n487_n553# a_487_n465# a_n29_n465# a_n679_n687# a_29_n553# a_n287_n465#
X0 a_487_n465# a_287_n553# a_229_n465# a_n679_n687# sky130_fd_pr__nfet_g5v0d10v5 ad=1.35 pd=9.88 as=0.674 ps=4.94 w=4.65 l=1
X1 a_229_n465# a_29_n553# a_n29_n465# a_n679_n687# sky130_fd_pr__nfet_g5v0d10v5 ad=0.674 pd=4.94 as=0.674 ps=4.94 w=4.65 l=1
X2 a_n29_n465# a_n229_n553# a_n287_n465# a_n679_n687# sky130_fd_pr__nfet_g5v0d10v5 ad=0.674 pd=4.94 as=0.674 ps=4.94 w=4.65 l=1
X3 a_n287_n465# a_n487_n553# a_n545_n465# a_n679_n687# sky130_fd_pr__nfet_g5v0d10v5 ad=0.674 pd=4.94 as=1.35 ps=9.88 w=4.65 l=1
C0 a_487_n465# a_287_n553# 0.105f
C1 a_n29_n465# a_n287_n465# 0.255f
C2 a_229_n465# a_287_n553# 0.105f
C3 a_29_n553# a_287_n553# 0.104f
C4 a_n487_n553# a_n287_n465# 0.105f
C5 a_n29_n465# a_n229_n553# 0.105f
C6 a_n545_n465# a_n287_n465# 0.255f
C7 a_n487_n553# a_n229_n553# 0.104f
C8 a_29_n553# a_n229_n553# 0.104f
C9 a_229_n465# a_n29_n465# 0.255f
C10 a_29_n553# a_n29_n465# 0.105f
C11 a_n487_n553# a_n545_n465# 0.105f
C12 a_229_n465# a_487_n465# 0.255f
C13 a_n229_n553# a_n287_n465# 0.105f
C14 a_229_n465# a_29_n553# 0.105f
C15 a_487_n465# a_n679_n687# 0.517f
C16 a_229_n465# a_n679_n687# 0.157f
C17 a_n29_n465# a_n679_n687# 0.157f
C18 a_n287_n465# a_n679_n687# 0.157f
C19 a_n545_n465# a_n679_n687# 0.517f
C20 a_287_n553# a_n679_n687# 0.651f
C21 a_29_n553# a_n679_n687# 0.588f
C22 a_n229_n553# a_n679_n687# 0.588f
C23 a_n487_n553# a_n679_n687# 0.651f
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_YPGNM4 a_545_n528# a_n545_n440# a_1577_n528#
+ a_1003_n440# a_n29_n440# a_29_n528# a_n1777_n528# a_487_n440# a_n745_n528# a_n1835_n440#
+ a_803_n528# a_n803_n440# a_1519_n440# a_1261_n440# a_n229_n528# a_n1319_n440# a_287_n528#
+ a_n1003_n528# a_n287_n440# a_n1061_n440# a_n1969_n662# a_745_n440# a_1319_n528#
+ a_1061_n528# a_1777_n440# a_n1519_n528# a_229_n440# a_n487_n528# a_n1261_n528# a_n1577_n440#
X0 a_1777_n440# a_1577_n528# a_1519_n440# a_n1969_n662# sky130_fd_pr__nfet_g5v0d10v5 ad=1.28 pd=9.38 as=0.638 ps=4.69 w=4.4 l=1
X1 a_1261_n440# a_1061_n528# a_1003_n440# a_n1969_n662# sky130_fd_pr__nfet_g5v0d10v5 ad=0.638 pd=4.69 as=0.638 ps=4.69 w=4.4 l=1
X2 a_229_n440# a_29_n528# a_n29_n440# a_n1969_n662# sky130_fd_pr__nfet_g5v0d10v5 ad=0.638 pd=4.69 as=0.638 ps=4.69 w=4.4 l=1
X3 a_n29_n440# a_n229_n528# a_n287_n440# a_n1969_n662# sky130_fd_pr__nfet_g5v0d10v5 ad=0.638 pd=4.69 as=0.638 ps=4.69 w=4.4 l=1
X4 a_n1319_n440# a_n1519_n528# a_n1577_n440# a_n1969_n662# sky130_fd_pr__nfet_g5v0d10v5 ad=0.638 pd=4.69 as=0.638 ps=4.69 w=4.4 l=1
X5 a_n545_n440# a_n745_n528# a_n803_n440# a_n1969_n662# sky130_fd_pr__nfet_g5v0d10v5 ad=0.638 pd=4.69 as=0.638 ps=4.69 w=4.4 l=1
X6 a_n803_n440# a_n1003_n528# a_n1061_n440# a_n1969_n662# sky130_fd_pr__nfet_g5v0d10v5 ad=0.638 pd=4.69 as=0.638 ps=4.69 w=4.4 l=1
X7 a_n287_n440# a_n487_n528# a_n545_n440# a_n1969_n662# sky130_fd_pr__nfet_g5v0d10v5 ad=0.638 pd=4.69 as=0.638 ps=4.69 w=4.4 l=1
X8 a_n1577_n440# a_n1777_n528# a_n1835_n440# a_n1969_n662# sky130_fd_pr__nfet_g5v0d10v5 ad=0.638 pd=4.69 as=1.28 ps=9.38 w=4.4 l=1
X9 a_1519_n440# a_1319_n528# a_1261_n440# a_n1969_n662# sky130_fd_pr__nfet_g5v0d10v5 ad=0.638 pd=4.69 as=0.638 ps=4.69 w=4.4 l=1
X10 a_n1061_n440# a_n1261_n528# a_n1319_n440# a_n1969_n662# sky130_fd_pr__nfet_g5v0d10v5 ad=0.638 pd=4.69 as=0.638 ps=4.69 w=4.4 l=1
X11 a_1003_n440# a_803_n528# a_745_n440# a_n1969_n662# sky130_fd_pr__nfet_g5v0d10v5 ad=0.638 pd=4.69 as=0.638 ps=4.69 w=4.4 l=1
X12 a_487_n440# a_287_n528# a_229_n440# a_n1969_n662# sky130_fd_pr__nfet_g5v0d10v5 ad=0.638 pd=4.69 as=0.638 ps=4.69 w=4.4 l=1
X13 a_745_n440# a_545_n528# a_487_n440# a_n1969_n662# sky130_fd_pr__nfet_g5v0d10v5 ad=0.638 pd=4.69 as=0.638 ps=4.69 w=4.4 l=1
C0 a_1519_n440# a_1261_n440# 0.241f
C1 a_745_n440# a_487_n440# 0.241f
C2 a_n745_n528# a_n1003_n528# 0.104f
C3 a_n803_n440# a_n1003_n528# 0.0995f
C4 a_n803_n440# a_n745_n528# 0.0995f
C5 a_n545_n440# a_n745_n528# 0.0995f
C6 a_1319_n528# a_1577_n528# 0.104f
C7 a_n803_n440# a_n545_n440# 0.241f
C8 a_803_n528# a_1061_n528# 0.104f
C9 a_287_n528# a_29_n528# 0.104f
C10 a_n229_n528# a_29_n528# 0.104f
C11 a_n1519_n528# a_n1319_n440# 0.0995f
C12 a_1319_n528# a_1519_n440# 0.0995f
C13 a_n229_n528# a_n287_n440# 0.0995f
C14 a_803_n528# a_1003_n440# 0.0995f
C15 a_n487_n528# a_n745_n528# 0.104f
C16 a_n1061_n440# a_n1003_n528# 0.0995f
C17 a_n545_n440# a_n487_n528# 0.0995f
C18 a_n1577_n440# a_n1519_n528# 0.0995f
C19 a_n803_n440# a_n1061_n440# 0.241f
C20 a_n1577_n440# a_n1777_n528# 0.0995f
C21 a_29_n528# a_n29_n440# 0.0995f
C22 a_n1577_n440# a_n1835_n440# 0.241f
C23 a_803_n528# a_545_n528# 0.104f
C24 a_n287_n440# a_n29_n440# 0.241f
C25 a_545_n528# a_487_n440# 0.0995f
C26 a_1319_n528# a_1261_n440# 0.0995f
C27 a_1061_n528# a_1261_n440# 0.0995f
C28 a_n1061_n440# a_n1319_n440# 0.241f
C29 a_n1261_n528# a_n1519_n528# 0.104f
C30 a_229_n440# a_487_n440# 0.241f
C31 a_n229_n528# a_n29_n440# 0.0995f
C32 a_1319_n528# a_1061_n528# 0.104f
C33 a_n1261_n528# a_n1003_n528# 0.104f
C34 a_n545_n440# a_n287_n440# 0.241f
C35 a_n1577_n440# a_n1319_n440# 0.241f
C36 a_229_n440# a_29_n528# 0.0995f
C37 a_1261_n440# a_1003_n440# 0.241f
C38 a_1519_n440# a_1577_n528# 0.0995f
C39 a_1003_n440# a_745_n440# 0.241f
C40 a_287_n528# a_545_n528# 0.104f
C41 a_1061_n528# a_1003_n440# 0.0995f
C42 a_229_n440# a_287_n528# 0.0995f
C43 a_745_n440# a_545_n528# 0.0995f
C44 a_n1261_n528# a_n1319_n440# 0.0995f
C45 a_n287_n440# a_n487_n528# 0.0995f
C46 a_n1777_n528# a_n1519_n528# 0.104f
C47 a_n1261_n528# a_n1061_n440# 0.0995f
C48 a_n229_n528# a_n487_n528# 0.104f
C49 a_n1777_n528# a_n1835_n440# 0.0995f
C50 a_1777_n440# a_1577_n528# 0.0995f
C51 a_1777_n440# a_1519_n440# 0.241f
C52 a_803_n528# a_745_n440# 0.0995f
C53 a_287_n528# a_487_n440# 0.0995f
C54 a_229_n440# a_n29_n440# 0.241f
C55 a_1777_n440# a_n1969_n662# 0.491f
C56 a_1519_n440# a_n1969_n662# 0.15f
C57 a_1261_n440# a_n1969_n662# 0.15f
C58 a_1003_n440# a_n1969_n662# 0.15f
C59 a_745_n440# a_n1969_n662# 0.15f
C60 a_487_n440# a_n1969_n662# 0.15f
C61 a_229_n440# a_n1969_n662# 0.15f
C62 a_n29_n440# a_n1969_n662# 0.15f
C63 a_n287_n440# a_n1969_n662# 0.15f
C64 a_n545_n440# a_n1969_n662# 0.15f
C65 a_n803_n440# a_n1969_n662# 0.15f
C66 a_n1061_n440# a_n1969_n662# 0.15f
C67 a_n1319_n440# a_n1969_n662# 0.15f
C68 a_n1577_n440# a_n1969_n662# 0.15f
C69 a_n1835_n440# a_n1969_n662# 0.491f
C70 a_1577_n528# a_n1969_n662# 0.65f
C71 a_1319_n528# a_n1969_n662# 0.587f
C72 a_1061_n528# a_n1969_n662# 0.587f
C73 a_803_n528# a_n1969_n662# 0.587f
C74 a_545_n528# a_n1969_n662# 0.587f
C75 a_287_n528# a_n1969_n662# 0.587f
C76 a_29_n528# a_n1969_n662# 0.587f
C77 a_n229_n528# a_n1969_n662# 0.587f
C78 a_n487_n528# a_n1969_n662# 0.587f
C79 a_n745_n528# a_n1969_n662# 0.587f
C80 a_n1003_n528# a_n1969_n662# 0.587f
C81 a_n1261_n528# a_n1969_n662# 0.587f
C82 a_n1519_n528# a_n1969_n662# 0.587f
C83 a_n1777_n528# a_n1969_n662# 0.65f
.ends

.subckt RB_array_20 VDD R1 D0 m1_2124_1470# m1_5470_410# m1_2651_1472# m1_3160_410#
+ m1_4060_410# D3 D1 R2 D4 D2 VSS m1_7940_410#
XXR1 VSS R2 m1_2651_1472# sky130_fd_pr__res_high_po_0p69_JKKHRG
XXR2 VSS R2 m1_2124_1470# sky130_fd_pr__res_high_po_0p69_JKKHRG
XXR3 R2 m1_3160_410# R2 VSS m1_3160_410# sky130_fd_pr__res_high_po_0p69_Z3RMRJ
XXR5 m1_5470_410# R2 R2 R2 m1_5470_410# R2 R2 m1_5470_410# R2 m1_5470_410# m1_5470_410#
+ m1_5470_410# m1_5470_410# R2 VSS R2 m1_5470_410# sky130_fd_pr__res_high_po_0p69_Z3RMR6
XXR4 R2 VSS m1_4060_410# R2 R2 m1_4060_410# m1_4060_410# m1_4060_410# R2 sky130_fd_pr__res_high_po_0p69_YMHKRJ
XXR6 m1_7940_410# R2 R2 R2 R2 m1_7940_410# m1_7940_410# m1_7940_410# R2 VSS R2 R2
+ m1_7940_410# R2 m1_7940_410# R2 R2 m1_7940_410# m1_7940_410# R2 R2 R2 m1_7940_410#
+ m1_7940_410# m1_7940_410# m1_7940_410# R2 R2 m1_7940_410# m1_7940_410# R2 m1_7940_410#
+ m1_7940_410# sky130_fd_pr__res_high_po_0p69_HBQF5Z
XXM6 D0 m1_2651_1472# VSS R1 sky130_fd_pr__nfet_g5v0d10v5_727CUP
XXM7 m1_3160_410# VSS D1 m1_3160_410# R1 D1 sky130_fd_pr__nfet_g5v0d10v5_VU5C5A
XXM9 m1_5470_410# R1 D3 D3 R1 m1_5470_410# D3 R1 D3 D3 D3 R1 m1_5470_410# m1_5470_410#
+ D3 VSS D3 m1_5470_410# sky130_fd_pr__nfet_g5v0d10v5_J97EKB
XXM8 D2 D2 R1 m1_4060_410# D2 m1_4060_410# m1_4060_410# VSS D2 R1 sky130_fd_pr__nfet_g5v0d10v5_S7E57E
XXM10 D4 R1 D4 R1 R1 D4 D4 R1 D4 m1_7940_410# D4 m1_7940_410# R1 m1_7940_410# D4 m1_7940_410#
+ D4 D4 m1_7940_410# R1 VSS m1_7940_410# D4 D4 m1_7940_410# D4 m1_7940_410# D4 D4
+ R1 sky130_fd_pr__nfet_g5v0d10v5_YPGNM4
XXM11 VDD m1_2124_1470# VSS R1 sky130_fd_pr__nfet_g5v0d10v5_727CUP
C0 D0 m1_4060_410# 7.28e-21
C1 D3 D0 0.0725f
C2 m1_2651_1472# m1_4060_410# 2.22e-21
C3 D3 m1_2651_1472# 0.0446f
C4 D3 VDD 0.0728f
C5 m1_5470_410# D4 1.37f
C6 D0 D2 0.0732f
C7 D4 m1_4060_410# 0.742f
C8 D3 D4 3.99f
C9 m1_2651_1472# D2 0.0483f
C10 D4 m1_7940_410# 8.65f
C11 VDD D2 0.0734f
C12 m1_5470_410# R1 0.379f
C13 R1 m1_4060_410# 0.226f
C14 D3 R1 4.08f
C15 m1_3160_410# m1_4060_410# 0.201f
C16 R1 m1_7940_410# 0.29f
C17 D4 D2 0.308f
C18 D3 m1_3160_410# 0.12f
C19 R1 D2 2.15f
C20 m1_3160_410# D2 0.163f
C21 D0 m1_2651_1472# 0.449f
C22 D0 VDD 0.332f
C23 D4 D0 0.0964f
C24 D3 m1_2124_1470# 0.0433f
C25 D4 m1_2651_1472# 0.0516f
C26 D4 VDD 0.0966f
C27 D1 m1_4060_410# 1.86e-19
C28 R1 D0 0.619f
C29 D3 D1 0.145f
C30 m1_3160_410# D0 0.00189f
C31 m1_2124_1470# D2 0.0469f
C32 R1 m1_2651_1472# -0.107f
C33 R1 VDD 0.551f
C34 m1_3160_410# m1_2651_1472# 0.19f
C35 m1_3160_410# VDD 4.48e-19
C36 D1 D2 1.31f
C37 R1 D4 7.57f
C38 m1_3160_410# D4 0.458f
C39 m1_3160_410# R1 0.177f
C40 D0 m1_2124_1470# 0.126f
C41 m1_2124_1470# m1_2651_1472# 0.104f
C42 m1_2124_1470# VDD 0.494f
C43 D1 D0 0.731f
C44 D1 m1_2651_1472# 0.114f
C45 D1 VDD 0.0754f
C46 D4 m1_2124_1470# 0.0503f
C47 D4 D1 0.154f
C48 R1 m1_2124_1470# 0.0621f
C49 m1_3160_410# m1_2124_1470# 1.43e-19
C50 R1 D1 1.16f
C51 m1_3160_410# D1 1.09f
C52 m1_5470_410# m1_4060_410# 0.176f
C53 D3 m1_5470_410# 3.93f
C54 m1_5470_410# m1_7940_410# 0.197f
C55 D3 m1_4060_410# 0.2f
C56 D3 m1_7940_410# 5.93e-19
C57 m1_5470_410# D2 5.82e-19
C58 D2 m1_4060_410# 2.08f
C59 D3 D2 2.27f
C60 D1 m1_2124_1470# 0.0674f
C61 R1 VSS 4.54f
C62 VDD VSS 0.914f
C63 m1_7940_410# VSS 7.18f
C64 D4 VSS 8.99f
C65 D2 VSS 2.7f
C66 D3 VSS 5.24f
C67 D1 VSS 1.48f
C68 D0 VSS 0.884f
C69 m1_4060_410# VSS 3.17f
C70 m1_5470_410# VSS 4.68f
C71 m1_3160_410# VSS 2.43f
C72 R2 VSS 15.3f
C73 m1_2124_1470# VSS 1.55f
C74 m1_2651_1472# VSS 1.58f
.ends

.subckt sky130_fd_pr__res_high_po_0p69_T8KQH6 a_n199_n866# a_n69_n736# a_n69_304#
X0 a_n69_304# a_n69_n736# a_n199_n866# sky130_fd_pr__res_high_po_0p69 l=3.04
C0 a_n69_n736# a_n69_304# 0.0134f
C1 a_n69_n736# a_n199_n866# 0.659f
C2 a_n69_304# a_n199_n866# 0.659f
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_K8DQNF a_n29_n1536# a_229_n1536# a_n229_n1562#
+ w_n487_n1762# a_n287_n1536# a_29_n1562# VSUBS
X0 a_n29_n1536# a_n229_n1562# a_n287_n1536# w_n487_n1762# sky130_fd_pr__pfet_g5v0d10v5 ad=2.17 pd=15.3 as=4.35 ps=30.6 w=15 l=1
X1 a_229_n1536# a_29_n1562# a_n29_n1536# w_n487_n1762# sky130_fd_pr__pfet_g5v0d10v5 ad=4.35 pd=30.6 as=2.17 ps=15.3 w=15 l=1
C0 a_29_n1562# w_n487_n1762# 0.257f
C1 a_n229_n1562# w_n487_n1762# 0.257f
C2 a_n29_n1536# a_n287_n1536# 0.82f
C3 w_n487_n1762# a_229_n1536# 0.868f
C4 a_n29_n1536# w_n487_n1762# 0.023f
C5 a_n229_n1562# a_29_n1562# 0.0619f
C6 a_29_n1562# a_229_n1536# 0.326f
C7 a_29_n1562# a_n29_n1536# 0.326f
C8 a_n229_n1562# a_n29_n1536# 0.326f
C9 a_n29_n1536# a_229_n1536# 0.82f
C10 a_n287_n1536# w_n487_n1762# 0.868f
C11 a_n229_n1562# a_n287_n1536# 0.326f
C12 a_229_n1536# VSUBS 0.733f
C13 a_n29_n1536# VSUBS 0.418f
C14 a_n287_n1536# VSUBS 0.733f
C15 a_29_n1562# VSUBS 0.228f
C16 a_n229_n1562# VSUBS 0.228f
C17 w_n487_n1762# VSUBS 12.4f
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_VYCZE8 a_100_n1681# a_n292_n1841# a_n100_n1707#
+ a_n158_n1681#
X0 a_100_n1681# a_n100_n1707# a_n158_n1681# a_n292_n1841# sky130_fd_pr__nfet_g5v0d10v5 ad=4.78 pd=33.6 as=4.78 ps=33.6 w=16.5 l=1
C0 a_100_n1681# a_n100_n1707# 0.358f
C1 a_n158_n1681# a_n100_n1707# 0.358f
C2 a_n158_n1681# a_100_n1681# 0.901f
C3 a_100_n1681# a_n292_n1841# 1.75f
C4 a_n158_n1681# a_n292_n1841# 1.75f
C5 a_n100_n1707# a_n292_n1841# 0.513f
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_F3SB2X a_n100_n1632# a_100_n1544# a_n292_n1766#
+ a_n158_n1544#
X0 a_100_n1544# a_n100_n1632# a_n158_n1544# a_n292_n1766# sky130_fd_pr__nfet_g5v0d10v5 ad=4.48 pd=31.5 as=4.48 ps=31.5 w=15.4 l=1
C0 a_100_n1544# a_n100_n1632# 0.335f
C1 a_n158_n1544# a_n100_n1632# 0.335f
C2 a_n158_n1544# a_100_n1544# 0.844f
C3 a_100_n1544# a_n292_n1766# 1.64f
C4 a_n158_n1544# a_n292_n1766# 1.64f
C5 a_n100_n1632# a_n292_n1766# 0.743f
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_2HXNYY a_n158_n1900# a_100_n1900# a_n292_n2122#
+ a_n100_n1988#
X0 a_100_n1900# a_n100_n1988# a_n158_n1900# a_n292_n2122# sky130_fd_pr__nfet_g5v0d10v5 ad=5.51 pd=38.6 as=5.51 ps=38.6 w=19 l=1
C0 a_100_n1900# a_n100_n1988# 0.411f
C1 a_n158_n1900# a_n100_n1988# 0.411f
C2 a_n158_n1900# a_100_n1900# 1.04f
C3 a_100_n1900# a_n292_n2122# 2.01f
C4 a_n158_n1900# a_n292_n2122# 2.01f
C5 a_n100_n1988# a_n292_n2122# 0.743f
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_24QKAW a_29_n1997# a_n487_n1997# a_487_n1900#
+ a_n287_n1900# a_n229_n1997# a_n545_n1900# a_n29_n1900# a_287_n1997# w_n745_n2197#
+ a_229_n1900# VSUBS
X0 a_487_n1900# a_287_n1997# a_229_n1900# w_n745_n2197# sky130_fd_pr__pfet_g5v0d10v5 ad=5.51 pd=38.6 as=2.76 ps=19.3 w=19 l=1
X1 a_n287_n1900# a_n487_n1997# a_n545_n1900# w_n745_n2197# sky130_fd_pr__pfet_g5v0d10v5 ad=2.76 pd=19.3 as=5.51 ps=38.6 w=19 l=1
X2 a_n29_n1900# a_n229_n1997# a_n287_n1900# w_n745_n2197# sky130_fd_pr__pfet_g5v0d10v5 ad=2.76 pd=19.3 as=2.76 ps=19.3 w=19 l=1
X3 a_229_n1900# a_29_n1997# a_n29_n1900# w_n745_n2197# sky130_fd_pr__pfet_g5v0d10v5 ad=2.76 pd=19.3 as=2.76 ps=19.3 w=19 l=1
C0 a_n229_n1997# a_n29_n1900# 0.411f
C1 a_n287_n1900# a_n229_n1997# 0.411f
C2 a_n287_n1900# a_n487_n1997# 0.411f
C3 a_n287_n1900# a_n545_n1900# 1.04f
C4 a_n229_n1997# w_n745_n2197# 0.343f
C5 a_n487_n1997# w_n745_n2197# 0.386f
C6 a_287_n1997# a_29_n1997# 0.109f
C7 w_n745_n2197# a_n545_n1900# 1.09f
C8 a_487_n1900# a_287_n1997# 0.411f
C9 a_287_n1997# w_n745_n2197# 0.386f
C10 a_n487_n1997# a_n229_n1997# 0.109f
C11 a_229_n1900# a_29_n1997# 0.411f
C12 a_n487_n1997# a_n545_n1900# 0.411f
C13 a_229_n1900# a_n29_n1900# 1.04f
C14 a_229_n1900# a_487_n1900# 1.04f
C15 a_229_n1900# w_n745_n2197# 0.022f
C16 a_29_n1997# a_n29_n1900# 0.411f
C17 a_229_n1900# a_287_n1997# 0.411f
C18 a_n287_n1900# a_n29_n1900# 1.04f
C19 a_29_n1997# w_n745_n2197# 0.343f
C20 a_n29_n1900# w_n745_n2197# 0.022f
C21 a_n287_n1900# w_n745_n2197# 0.022f
C22 a_487_n1900# w_n745_n2197# 1.09f
C23 a_n229_n1997# a_29_n1997# 0.109f
C24 a_487_n1900# VSUBS 0.925f
C25 a_229_n1900# VSUBS 0.527f
C26 a_n29_n1900# VSUBS 0.527f
C27 a_n287_n1900# VSUBS 0.527f
C28 a_n545_n1900# VSUBS 0.925f
C29 a_287_n1997# VSUBS 0.311f
C30 a_29_n1997# VSUBS 0.288f
C31 a_n229_n1997# VSUBS 0.288f
C32 a_n487_n1997# VSUBS 0.311f
C33 w_n745_n2197# VSUBS 22.5f
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_LB7Y8R a_n100_n157# a_n158_n69# a_n292_n291#
+ a_100_n69#
X0 a_100_n69# a_n100_n157# a_n158_n69# a_n292_n291# sky130_fd_pr__nfet_g5v0d10v5 ad=0.2 pd=1.96 as=0.2 ps=1.96 w=0.69 l=1
C0 a_100_n69# a_n100_n157# 0.0202f
C1 a_n100_n157# a_n158_n69# 0.0202f
C2 a_100_n69# a_n158_n69# 0.0387f
C3 a_100_n69# a_n292_n291# 0.105f
C4 a_n158_n69# a_n292_n291# 0.105f
C5 a_n100_n157# a_n292_n291# 0.683f
.ends

.subckt sky130_fd_pr__cap_mim_m3_1_8DB3RK m3_n876_n730# c1_n836_n690# VSUBS
X0 c1_n836_n690# m3_n876_n730# sky130_fd_pr__cap_mim_m3_1 l=6.9 w=6.9
C0 m3_n876_n730# c1_n836_n690# 4.73f
C1 c1_n836_n690# VSUBS 0.686f
C2 m3_n876_n730# VSUBS 2.42f
.ends

.subckt opamp V2 VOUT a_4864_8007# V1 m1_4128_540# VDD m1_5284_1188# m1_4306_994#
+ m3_5211_1261# VSS m1_5053_7611#
XXR3 VSS m1_4128_540# VOUT sky130_fd_pr__res_high_po_0p69_T8KQH6
XXM1 m1_5053_7611# VDD a_4864_8007# VDD VDD a_4864_8007# VSS sky130_fd_pr__pfet_g5v0d10v5_K8DQNF
XXM2 m1_4306_994# VSS V2 a_4864_8007# sky130_fd_pr__nfet_g5v0d10v5_VYCZE8
XXM3 a_4864_8007# VDD a_4864_8007# VDD VDD a_4864_8007# VSS sky130_fd_pr__pfet_g5v0d10v5_K8DQNF
XXM4 m1_5053_7611# VSS V1 m1_4306_994# sky130_fd_pr__nfet_g5v0d10v5_VYCZE8
XXM5 m1_5284_1188# VSS VSS m1_4306_994# sky130_fd_pr__nfet_g5v0d10v5_F3SB2X
XXM6 VSS VOUT VSS m1_5284_1188# sky130_fd_pr__nfet_g5v0d10v5_2HXNYY
XXM7 m1_5284_1188# m1_5284_1188# VSS VSS sky130_fd_pr__nfet_g5v0d10v5_F3SB2X
XXM8 m1_5053_7611# m1_5053_7611# VDD VOUT m1_5053_7611# VDD VDD m1_5053_7611# VDD
+ VOUT VSS sky130_fd_pr__pfet_g5v0d10v5_24QKAW
XXM9 VDD VDD VSS m1_5284_1188# sky130_fd_pr__nfet_g5v0d10v5_LB7Y8R
XXC1 m1_5053_7611# m1_4128_540# VSS sky130_fd_pr__cap_mim_m3_1_8DB3RK
C0 V2 V1 0.16f
C1 m1_5284_1188# V1 0.00363f
C2 a_4864_8007# V2 0.263f
C3 a_4864_8007# m1_5284_1188# 0.00623f
C4 m1_5053_7611# V2 4.01e-19
C5 m1_5284_1188# m1_5053_7611# 0.0361f
C6 m3_5211_1261# m1_4306_994# 0.771f
C7 m1_4128_540# V2 0.179f
C8 m1_4128_540# m1_5284_1188# 0.031f
C9 VDD V2 0.00314f
C10 m1_5284_1188# VDD 1.67f
C11 VOUT m1_5284_1188# 2.28f
C12 a_4864_8007# V1 0.283f
C13 m1_5053_7611# V1 0.143f
C14 m1_4128_540# V1 0.088f
C15 a_4864_8007# m1_5053_7611# 1.78f
C16 VDD V1 0.275f
C17 m1_4306_994# V2 0.213f
C18 m1_5284_1188# m1_4306_994# 2.09f
C19 m3_5211_1261# V2 0.0767f
C20 m3_5211_1261# m1_5284_1188# 0.446f
C21 a_4864_8007# m1_4128_540# 0.503f
C22 VOUT V1 2.75e-19
C23 m1_4128_540# m1_5053_7611# 0.115f
C24 a_4864_8007# VDD 1.96f
C25 VDD m1_5053_7611# 10.4f
C26 a_4864_8007# VOUT 0.00842f
C27 VOUT m1_5053_7611# 7.29f
C28 m1_4128_540# VDD 0.376f
C29 VOUT m1_4128_540# 0.00888f
C30 m1_4306_994# V1 0.399f
C31 m3_5211_1261# V1 0.14f
C32 VOUT VDD -1.29f
C33 a_4864_8007# m1_4306_994# 0.127f
C34 a_4864_8007# m3_5211_1261# 0.0192f
C35 m1_5284_1188# V2 9.56e-20
C36 m1_5053_7611# m1_4306_994# 0.673f
C37 m3_5211_1261# m1_5053_7611# 0.0415f
C38 m1_4128_540# m1_4306_994# 0.354f
C39 m3_5211_1261# m1_4128_540# 0.0111f
C40 VDD m1_4306_994# 0.00701f
C41 m3_5211_1261# VDD 0.0192f
C42 VOUT m1_4306_994# 0.00433f
C43 m3_5211_1261# VOUT 0.00865f
C44 m3_5211_1261# VSS 1.23f
C45 VDD VSS 46.6f
C46 m1_5053_7611# VSS 4.65f
C47 VOUT VSS 4.32f
C48 m1_5284_1188# VSS 8.17f
C49 V1 VSS 0.865f
C50 m1_4306_994# VSS 5.55f
C51 V2 VSS 0.848f
C52 a_4864_8007# VSS 4.88f
C53 m1_4128_540# VSS 2.47f
.ends

.subckt sky130_fd_pr__res_high_po_0p69_WX3C5M a_2856_n1638# a_3090_1206# a_n3930_1206#
+ a_n5100_n1638# a_4260_n1638# a_7068_1206# a_516_n1638# a_6600_1206# a_n654_1206#
+ a_48_1206# a_4728_n1638# a_5196_1206# a_6132_n1638# a_n2526_1206# a_n6972_n1638#
+ a_5430_n1638# a_n5100_1206# a_3324_1206# a_6834_1206# a_7302_n1638# a_6600_n1638#
+ a_n888_1206# a_n7206_1206# a_n1122_n1638# a_1452_1206# a_4962_1206# a_n5334_1206#
+ a_n4398_n1638# a_n186_n1638# a_n3696_n1638# a_n2994_n1638# a_2154_n1638# a_n3462_1206#
+ a_n6972_1206# a_1452_n1638# a_3558_1206# a_6132_1206# a_n186_1206# a_n5568_n1638#
+ a_n1590_1206# a_n4866_n1638# a_1686_1206# a_4026_n1638# a_750_1206# a_3324_n1638#
+ a_n654_n1638# a_n2058_1206# a_n5568_1206# a_n6270_n1638# a_4260_1206# a_2622_n1638#
+ a_1920_n1638# a_984_n1638# a_n6738_n1638# a_n3696_1206# a_5898_n1638# a_n6270_1206#
+ a_6366_1206# a_n7440_n1638# a_984_1206# a_4494_1206# a_n1824_1206# a_n2292_n1638#
+ a_n1590_n1638# a_2622_1206# a_n6504_1206# a_1218_n1638# a_282_1206# a_n4164_n1638#
+ a_n3462_n1638# a_n2760_n1638# a_n1122_1206# a_n4632_1206# a_282_n1638# a_1218_1206#
+ a_4728_1206# a_7302_1206# a_n6036_n1638# a_5196_n1638# a_n5334_n1638# a_48_n1638#
+ a_n2760_1206# a_2856_1206# a_4494_n1638# a_n4632_n1638# a_3792_n1638# a_n3228_1206#
+ a_n3930_n1638# a_n6738_1206# a_n420_n1638# a_5430_1206# a_750_n1638# a_7068_n1638#
+ a_n7206_n1638# a_6366_n1638# a_n1356_1206# a_n4866_1206# a_n6504_n1638# a_5664_n1638#
+ a_n5802_n1638# a_516_1206# a_n7440_1206# a_4962_n1638# a_4026_1206# a_n7570_n1768#
+ a_n2994_1206# a_2154_1206# a_5664_1206# a_6834_n1638# a_n6036_1206# a_n2058_n1638#
+ a_n1356_n1638# a_3792_1206# a_n4164_1206# a_n3228_n1638# a_2388_n1638# a_n2526_n1638#
+ a_n420_1206# a_n2292_1206# a_1686_n1638# a_2388_1206# a_5898_1206# a_n1824_n1638#
+ a_3090_n1638# a_1920_1206# a_n5802_1206# a_3558_n1638# a_n888_n1638# a_n4398_1206#
X0 a_n420_1206# a_n420_n1638# a_n7570_n1768# sky130_fd_pr__res_high_po_0p69 l=12.1
X1 a_3090_1206# a_3090_n1638# a_n7570_n1768# sky130_fd_pr__res_high_po_0p69 l=12.1
X2 a_n6036_1206# a_n6036_n1638# a_n7570_n1768# sky130_fd_pr__res_high_po_0p69 l=12.1
X3 a_n2058_1206# a_n2058_n1638# a_n7570_n1768# sky130_fd_pr__res_high_po_0p69 l=12.1
X4 a_1452_1206# a_1452_n1638# a_n7570_n1768# sky130_fd_pr__res_high_po_0p69 l=12.1
X5 a_5430_1206# a_5430_n1638# a_n7570_n1768# sky130_fd_pr__res_high_po_0p69 l=12.1
X6 a_5196_1206# a_5196_n1638# a_n7570_n1768# sky130_fd_pr__res_high_po_0p69 l=12.1
X7 a_n3696_1206# a_n3696_n1638# a_n7570_n1768# sky130_fd_pr__res_high_po_0p69 l=12.1
X8 a_3558_1206# a_3558_n1638# a_n7570_n1768# sky130_fd_pr__res_high_po_0p69 l=12.1
X9 a_n3462_1206# a_n3462_n1638# a_n7570_n1768# sky130_fd_pr__res_high_po_0p69 l=12.1
X10 a_3324_1206# a_3324_n1638# a_n7570_n1768# sky130_fd_pr__res_high_po_0p69 l=12.1
X11 a_7068_1206# a_7068_n1638# a_n7570_n1768# sky130_fd_pr__res_high_po_0p69 l=12.1
X12 a_7302_1206# a_7302_n1638# a_n7570_n1768# sky130_fd_pr__res_high_po_0p69 l=12.1
X13 a_n5802_1206# a_n5802_n1638# a_n7570_n1768# sky130_fd_pr__res_high_po_0p69 l=12.1
X14 a_n1824_1206# a_n1824_n1638# a_n7570_n1768# sky130_fd_pr__res_high_po_0p69 l=12.1
X15 a_n5568_1206# a_n5568_n1638# a_n7570_n1768# sky130_fd_pr__res_high_po_0p69 l=12.1
X16 a_n1590_1206# a_n1590_n1638# a_n7570_n1768# sky130_fd_pr__res_high_po_0p69 l=12.1
X17 a_4962_1206# a_4962_n1638# a_n7570_n1768# sky130_fd_pr__res_high_po_0p69 l=12.1
X18 a_48_1206# a_48_n1638# a_n7570_n1768# sky130_fd_pr__res_high_po_0p69 l=12.1
X19 a_n3930_1206# a_n3930_n1638# a_n7570_n1768# sky130_fd_pr__res_high_po_0p69 l=12.1
X20 a_984_1206# a_984_n1638# a_n7570_n1768# sky130_fd_pr__res_high_po_0p69 l=12.1
X21 a_n5334_1206# a_n5334_n1638# a_n7570_n1768# sky130_fd_pr__res_high_po_0p69 l=12.1
X22 a_n1356_1206# a_n1356_n1638# a_n7570_n1768# sky130_fd_pr__res_high_po_0p69 l=12.1
X23 a_n5100_1206# a_n5100_n1638# a_n7570_n1768# sky130_fd_pr__res_high_po_0p69 l=12.1
X24 a_1218_1206# a_1218_n1638# a_n7570_n1768# sky130_fd_pr__res_high_po_0p69 l=12.1
X25 a_4494_1206# a_4494_n1638# a_n7570_n1768# sky130_fd_pr__res_high_po_0p69 l=12.1
X26 a_n6972_1206# a_n6972_n1638# a_n7570_n1768# sky130_fd_pr__res_high_po_0p69 l=12.1
X27 a_n2994_1206# a_n2994_n1638# a_n7570_n1768# sky130_fd_pr__res_high_po_0p69 l=12.1
X28 a_6834_1206# a_6834_n1638# a_n7570_n1768# sky130_fd_pr__res_high_po_0p69 l=12.1
X29 a_n7440_1206# a_n7440_n1638# a_n7570_n1768# sky130_fd_pr__res_high_po_0p69 l=12.1
X30 a_750_1206# a_750_n1638# a_n7570_n1768# sky130_fd_pr__res_high_po_0p69 l=12.1
X31 a_2856_1206# a_2856_n1638# a_n7570_n1768# sky130_fd_pr__res_high_po_0p69 l=12.1
X32 a_n1122_1206# a_n1122_n1638# a_n7570_n1768# sky130_fd_pr__res_high_po_0p69 l=12.1
X33 a_4260_1206# a_4260_n1638# a_n7570_n1768# sky130_fd_pr__res_high_po_0p69 l=12.1
X34 a_n888_1206# a_n888_n1638# a_n7570_n1768# sky130_fd_pr__res_high_po_0p69 l=12.1
X35 a_n7206_1206# a_n7206_n1638# a_n7570_n1768# sky130_fd_pr__res_high_po_0p69 l=12.1
X36 a_n3228_1206# a_n3228_n1638# a_n7570_n1768# sky130_fd_pr__res_high_po_0p69 l=12.1
X37 a_2622_1206# a_2622_n1638# a_n7570_n1768# sky130_fd_pr__res_high_po_0p69 l=12.1
X38 a_6366_1206# a_6366_n1638# a_n7570_n1768# sky130_fd_pr__res_high_po_0p69 l=12.1
X39 a_6600_1206# a_6600_n1638# a_n7570_n1768# sky130_fd_pr__res_high_po_0p69 l=12.1
X40 a_282_1206# a_282_n1638# a_n7570_n1768# sky130_fd_pr__res_high_po_0p69 l=12.1
X41 a_2388_1206# a_2388_n1638# a_n7570_n1768# sky130_fd_pr__res_high_po_0p69 l=12.1
X42 a_n4866_1206# a_n4866_n1638# a_n7570_n1768# sky130_fd_pr__res_high_po_0p69 l=12.1
X43 a_4728_1206# a_4728_n1638# a_n7570_n1768# sky130_fd_pr__res_high_po_0p69 l=12.1
X44 a_n654_1206# a_n654_n1638# a_n7570_n1768# sky130_fd_pr__res_high_po_0p69 l=12.1
X45 a_n2292_1206# a_n2292_n1638# a_n7570_n1768# sky130_fd_pr__res_high_po_0p69 l=12.1
X46 a_2154_1206# a_2154_n1638# a_n7570_n1768# sky130_fd_pr__res_high_po_0p69 l=12.1
X47 a_6132_1206# a_6132_n1638# a_n7570_n1768# sky130_fd_pr__res_high_po_0p69 l=12.1
X48 a_n4632_1206# a_n4632_n1638# a_n7570_n1768# sky130_fd_pr__res_high_po_0p69 l=12.1
X49 a_n4398_1206# a_n4398_n1638# a_n7570_n1768# sky130_fd_pr__res_high_po_0p69 l=12.1
X50 a_3792_1206# a_3792_n1638# a_n7570_n1768# sky130_fd_pr__res_high_po_0p69 l=12.1
X51 a_n186_1206# a_n186_n1638# a_n7570_n1768# sky130_fd_pr__res_high_po_0p69 l=12.1
X52 a_n6738_1206# a_n6738_n1638# a_n7570_n1768# sky130_fd_pr__res_high_po_0p69 l=12.1
X53 a_n2760_1206# a_n2760_n1638# a_n7570_n1768# sky130_fd_pr__res_high_po_0p69 l=12.1
X54 a_516_1206# a_516_n1638# a_n7570_n1768# sky130_fd_pr__res_high_po_0p69 l=12.1
X55 a_5898_1206# a_5898_n1638# a_n7570_n1768# sky130_fd_pr__res_high_po_0p69 l=12.1
X56 a_n4164_1206# a_n4164_n1638# a_n7570_n1768# sky130_fd_pr__res_high_po_0p69 l=12.1
X57 a_4026_1206# a_4026_n1638# a_n7570_n1768# sky130_fd_pr__res_high_po_0p69 l=12.1
X58 a_n6504_1206# a_n6504_n1638# a_n7570_n1768# sky130_fd_pr__res_high_po_0p69 l=12.1
X59 a_n2526_1206# a_n2526_n1638# a_n7570_n1768# sky130_fd_pr__res_high_po_0p69 l=12.1
X60 a_1920_1206# a_1920_n1638# a_n7570_n1768# sky130_fd_pr__res_high_po_0p69 l=12.1
X61 a_n6270_1206# a_n6270_n1638# a_n7570_n1768# sky130_fd_pr__res_high_po_0p69 l=12.1
X62 a_1686_1206# a_1686_n1638# a_n7570_n1768# sky130_fd_pr__res_high_po_0p69 l=12.1
X63 a_5664_1206# a_5664_n1638# a_n7570_n1768# sky130_fd_pr__res_high_po_0p69 l=12.1
C0 a_n6972_n1638# a_n6738_n1638# 0.296f
C1 a_n2760_n1638# a_n2526_n1638# 0.296f
C2 a_n5568_n1638# a_n5334_n1638# 0.296f
C3 a_516_1206# a_750_1206# 0.296f
C4 a_4026_1206# a_3792_1206# 0.296f
C5 a_2856_n1638# a_2622_n1638# 0.296f
C6 a_5898_n1638# a_5664_n1638# 0.296f
C7 a_n6036_1206# a_n5802_1206# 0.296f
C8 a_n6270_1206# a_n6504_1206# 0.296f
C9 a_48_1206# a_282_1206# 0.296f
C10 a_n5334_1206# a_n5568_1206# 0.296f
C11 a_4026_1206# a_4260_1206# 0.296f
C12 a_1920_1206# a_2154_1206# 0.296f
C13 a_4728_n1638# a_4494_n1638# 0.296f
C14 a_n2292_1206# a_n2526_1206# 0.296f
C15 a_n4632_n1638# a_n4866_n1638# 0.296f
C16 a_n1356_n1638# a_n1590_n1638# 0.296f
C17 a_1452_n1638# a_1686_n1638# 0.296f
C18 a_n4164_1206# a_n4398_1206# 0.296f
C19 a_n3462_1206# a_n3696_1206# 0.296f
C20 a_n6270_n1638# a_n6036_n1638# 0.296f
C21 a_5898_n1638# a_6132_n1638# 0.296f
C22 a_n3228_n1638# a_n2994_n1638# 0.296f
C23 a_3558_1206# a_3324_1206# 0.296f
C24 a_2856_1206# a_2622_1206# 0.296f
C25 a_6366_n1638# a_6600_n1638# 0.296f
C26 a_n1590_1206# a_n1824_1206# 0.296f
C27 a_n6036_1206# a_n6270_1206# 0.296f
C28 a_n3228_n1638# a_n3462_n1638# 0.296f
C29 a_6366_1206# a_6600_1206# 0.296f
C30 a_7302_n1638# a_7068_n1638# 0.296f
C31 a_n4632_1206# a_n4866_1206# 0.296f
C32 a_4026_n1638# a_3792_n1638# 0.296f
C33 a_n888_1206# a_n654_1206# 0.296f
C34 a_1218_1206# a_1452_1206# 0.296f
C35 a_n5100_n1638# a_n5334_n1638# 0.296f
C36 a_n1356_1206# a_n1122_1206# 0.296f
C37 a_4962_1206# a_5196_1206# 0.296f
C38 a_n1122_n1638# a_n888_n1638# 0.296f
C39 a_5430_n1638# a_5196_n1638# 0.296f
C40 a_n5100_n1638# a_n4866_n1638# 0.296f
C41 a_n2058_1206# a_n2292_1206# 0.296f
C42 a_n186_n1638# a_48_n1638# 0.296f
C43 a_6600_1206# a_6834_1206# 0.296f
C44 a_n420_1206# a_n654_1206# 0.296f
C45 a_n1122_n1638# a_n1356_n1638# 0.296f
C46 a_5430_n1638# a_5664_n1638# 0.296f
C47 a_n2760_n1638# a_n2994_n1638# 0.296f
C48 a_516_n1638# a_750_n1638# 0.296f
C49 a_2388_n1638# a_2622_n1638# 0.296f
C50 a_5664_1206# a_5430_1206# 0.296f
C51 a_1452_1206# a_1686_1206# 0.296f
C52 a_2154_1206# a_2388_1206# 0.296f
C53 a_n2058_n1638# a_n2292_n1638# 0.296f
C54 a_6366_1206# a_6132_1206# 0.296f
C55 a_4026_n1638# a_4260_n1638# 0.296f
C56 a_4260_1206# a_4494_1206# 0.296f
C57 a_48_n1638# a_282_n1638# 0.296f
C58 a_n1590_1206# a_n1356_1206# 0.296f
C59 a_984_n1638# a_1218_n1638# 0.296f
C60 a_3558_n1638# a_3324_n1638# 0.296f
C61 a_n186_n1638# a_n420_n1638# 0.296f
C62 a_1920_n1638# a_2154_n1638# 0.296f
C63 a_6834_n1638# a_6600_n1638# 0.296f
C64 a_6834_n1638# a_7068_n1638# 0.296f
C65 a_n6738_1206# a_n6972_1206# 0.296f
C66 a_n3930_n1638# a_n4164_n1638# 0.296f
C67 a_7068_1206# a_6834_1206# 0.296f
C68 a_n5568_1206# a_n5802_1206# 0.296f
C69 a_984_n1638# a_750_n1638# 0.296f
C70 a_n654_n1638# a_n420_n1638# 0.296f
C71 a_3792_1206# a_3558_1206# 0.296f
C72 a_2622_1206# a_2388_1206# 0.296f
C73 a_n3228_1206# a_n2994_1206# 0.296f
C74 a_n186_1206# a_48_1206# 0.296f
C75 a_n6738_1206# a_n6504_1206# 0.296f
C76 a_n2058_n1638# a_n1824_n1638# 0.296f
C77 a_n2058_1206# a_n1824_1206# 0.296f
C78 a_n6972_n1638# a_n7206_n1638# 0.296f
C79 a_n7206_1206# a_n6972_1206# 0.296f
C80 a_4962_n1638# a_5196_n1638# 0.296f
C81 a_1452_n1638# a_1218_n1638# 0.296f
C82 a_n2526_n1638# a_n2292_n1638# 0.296f
C83 a_516_1206# a_282_1206# 0.296f
C84 a_n5100_1206# a_n4866_1206# 0.296f
C85 a_4260_n1638# a_4494_n1638# 0.296f
C86 a_n888_n1638# a_n654_n1638# 0.296f
C87 a_1920_n1638# a_1686_n1638# 0.296f
C88 a_n3228_1206# a_n3462_1206# 0.296f
C89 a_3792_n1638# a_3558_n1638# 0.296f
C90 a_5898_1206# a_6132_1206# 0.296f
C91 a_3090_n1638# a_2856_n1638# 0.296f
C92 a_4962_n1638# a_4728_n1638# 0.296f
C93 a_n2760_1206# a_n2526_1206# 0.296f
C94 a_n5802_n1638# a_n6036_n1638# 0.296f
C95 a_n888_1206# a_n1122_1206# 0.296f
C96 a_5430_1206# a_5196_1206# 0.296f
C97 a_n7206_1206# a_n7440_1206# 0.296f
C98 a_n1590_n1638# a_n1824_n1638# 0.296f
C99 a_1218_1206# a_984_1206# 0.296f
C100 a_6366_n1638# a_6132_n1638# 0.296f
C101 a_n6270_n1638# a_n6504_n1638# 0.296f
C102 a_n5100_1206# a_n5334_1206# 0.296f
C103 a_3090_1206# a_3324_1206# 0.296f
C104 a_n3930_1206# a_n3696_1206# 0.296f
C105 a_n4632_n1638# a_n4398_n1638# 0.296f
C106 a_n3930_n1638# a_n3696_n1638# 0.296f
C107 a_984_1206# a_750_1206# 0.296f
C108 a_n2760_1206# a_n2994_1206# 0.296f
C109 a_n7206_n1638# a_n7440_n1638# 0.296f
C110 a_4728_1206# a_4494_1206# 0.296f
C111 a_n4164_n1638# a_n4398_n1638# 0.296f
C112 a_n3696_n1638# a_n3462_n1638# 0.296f
C113 a_n5568_n1638# a_n5802_n1638# 0.296f
C114 a_7068_1206# a_7302_1206# 0.296f
C115 a_3090_n1638# a_3324_n1638# 0.296f
C116 a_4962_1206# a_4728_1206# 0.296f
C117 a_1920_1206# a_1686_1206# 0.296f
C118 a_2388_n1638# a_2154_n1638# 0.296f
C119 a_n4632_1206# a_n4398_1206# 0.296f
C120 a_n186_1206# a_n420_1206# 0.296f
C121 a_3090_1206# a_2856_1206# 0.296f
C122 a_n4164_1206# a_n3930_1206# 0.296f
C123 a_516_n1638# a_282_n1638# 0.296f
C124 a_n6738_n1638# a_n6504_n1638# 0.296f
C125 a_5898_1206# a_5664_1206# 0.296f
C126 a_7302_n1638# a_n7570_n1768# 0.465f
C127 a_7302_1206# a_n7570_n1768# 0.465f
C128 a_7068_n1638# a_n7570_n1768# 0.255f
C129 a_7068_1206# a_n7570_n1768# 0.255f
C130 a_6834_n1638# a_n7570_n1768# 0.255f
C131 a_6834_1206# a_n7570_n1768# 0.255f
C132 a_6600_n1638# a_n7570_n1768# 0.255f
C133 a_6600_1206# a_n7570_n1768# 0.255f
C134 a_6366_n1638# a_n7570_n1768# 0.255f
C135 a_6366_1206# a_n7570_n1768# 0.255f
C136 a_6132_n1638# a_n7570_n1768# 0.255f
C137 a_6132_1206# a_n7570_n1768# 0.255f
C138 a_5898_n1638# a_n7570_n1768# 0.255f
C139 a_5898_1206# a_n7570_n1768# 0.255f
C140 a_5664_n1638# a_n7570_n1768# 0.255f
C141 a_5664_1206# a_n7570_n1768# 0.255f
C142 a_5430_n1638# a_n7570_n1768# 0.255f
C143 a_5430_1206# a_n7570_n1768# 0.255f
C144 a_5196_n1638# a_n7570_n1768# 0.255f
C145 a_5196_1206# a_n7570_n1768# 0.255f
C146 a_4962_n1638# a_n7570_n1768# 0.255f
C147 a_4962_1206# a_n7570_n1768# 0.255f
C148 a_4728_n1638# a_n7570_n1768# 0.255f
C149 a_4728_1206# a_n7570_n1768# 0.255f
C150 a_4494_n1638# a_n7570_n1768# 0.255f
C151 a_4494_1206# a_n7570_n1768# 0.255f
C152 a_4260_n1638# a_n7570_n1768# 0.255f
C153 a_4260_1206# a_n7570_n1768# 0.255f
C154 a_4026_n1638# a_n7570_n1768# 0.255f
C155 a_4026_1206# a_n7570_n1768# 0.255f
C156 a_3792_n1638# a_n7570_n1768# 0.255f
C157 a_3792_1206# a_n7570_n1768# 0.255f
C158 a_3558_n1638# a_n7570_n1768# 0.255f
C159 a_3558_1206# a_n7570_n1768# 0.255f
C160 a_3324_n1638# a_n7570_n1768# 0.255f
C161 a_3324_1206# a_n7570_n1768# 0.255f
C162 a_3090_n1638# a_n7570_n1768# 0.255f
C163 a_3090_1206# a_n7570_n1768# 0.255f
C164 a_2856_n1638# a_n7570_n1768# 0.255f
C165 a_2856_1206# a_n7570_n1768# 0.255f
C166 a_2622_n1638# a_n7570_n1768# 0.255f
C167 a_2622_1206# a_n7570_n1768# 0.255f
C168 a_2388_n1638# a_n7570_n1768# 0.255f
C169 a_2388_1206# a_n7570_n1768# 0.255f
C170 a_2154_n1638# a_n7570_n1768# 0.255f
C171 a_2154_1206# a_n7570_n1768# 0.255f
C172 a_1920_n1638# a_n7570_n1768# 0.255f
C173 a_1920_1206# a_n7570_n1768# 0.255f
C174 a_1686_n1638# a_n7570_n1768# 0.255f
C175 a_1686_1206# a_n7570_n1768# 0.255f
C176 a_1452_n1638# a_n7570_n1768# 0.255f
C177 a_1452_1206# a_n7570_n1768# 0.255f
C178 a_1218_n1638# a_n7570_n1768# 0.255f
C179 a_1218_1206# a_n7570_n1768# 0.255f
C180 a_984_n1638# a_n7570_n1768# 0.255f
C181 a_984_1206# a_n7570_n1768# 0.255f
C182 a_750_n1638# a_n7570_n1768# 0.255f
C183 a_750_1206# a_n7570_n1768# 0.255f
C184 a_516_n1638# a_n7570_n1768# 0.255f
C185 a_516_1206# a_n7570_n1768# 0.255f
C186 a_282_n1638# a_n7570_n1768# 0.255f
C187 a_282_1206# a_n7570_n1768# 0.255f
C188 a_48_n1638# a_n7570_n1768# 0.255f
C189 a_48_1206# a_n7570_n1768# 0.255f
C190 a_n186_n1638# a_n7570_n1768# 0.255f
C191 a_n186_1206# a_n7570_n1768# 0.255f
C192 a_n420_n1638# a_n7570_n1768# 0.255f
C193 a_n420_1206# a_n7570_n1768# 0.255f
C194 a_n654_n1638# a_n7570_n1768# 0.255f
C195 a_n654_1206# a_n7570_n1768# 0.255f
C196 a_n888_n1638# a_n7570_n1768# 0.255f
C197 a_n888_1206# a_n7570_n1768# 0.255f
C198 a_n1122_n1638# a_n7570_n1768# 0.255f
C199 a_n1122_1206# a_n7570_n1768# 0.255f
C200 a_n1356_n1638# a_n7570_n1768# 0.255f
C201 a_n1356_1206# a_n7570_n1768# 0.255f
C202 a_n1590_n1638# a_n7570_n1768# 0.255f
C203 a_n1590_1206# a_n7570_n1768# 0.255f
C204 a_n1824_n1638# a_n7570_n1768# 0.255f
C205 a_n1824_1206# a_n7570_n1768# 0.255f
C206 a_n2058_n1638# a_n7570_n1768# 0.255f
C207 a_n2058_1206# a_n7570_n1768# 0.255f
C208 a_n2292_n1638# a_n7570_n1768# 0.255f
C209 a_n2292_1206# a_n7570_n1768# 0.255f
C210 a_n2526_n1638# a_n7570_n1768# 0.255f
C211 a_n2526_1206# a_n7570_n1768# 0.255f
C212 a_n2760_n1638# a_n7570_n1768# 0.255f
C213 a_n2760_1206# a_n7570_n1768# 0.255f
C214 a_n2994_n1638# a_n7570_n1768# 0.255f
C215 a_n2994_1206# a_n7570_n1768# 0.255f
C216 a_n3228_n1638# a_n7570_n1768# 0.255f
C217 a_n3228_1206# a_n7570_n1768# 0.255f
C218 a_n3462_n1638# a_n7570_n1768# 0.255f
C219 a_n3462_1206# a_n7570_n1768# 0.255f
C220 a_n3696_n1638# a_n7570_n1768# 0.255f
C221 a_n3696_1206# a_n7570_n1768# 0.255f
C222 a_n3930_n1638# a_n7570_n1768# 0.255f
C223 a_n3930_1206# a_n7570_n1768# 0.255f
C224 a_n4164_n1638# a_n7570_n1768# 0.255f
C225 a_n4164_1206# a_n7570_n1768# 0.255f
C226 a_n4398_n1638# a_n7570_n1768# 0.255f
C227 a_n4398_1206# a_n7570_n1768# 0.255f
C228 a_n4632_n1638# a_n7570_n1768# 0.255f
C229 a_n4632_1206# a_n7570_n1768# 0.255f
C230 a_n4866_n1638# a_n7570_n1768# 0.255f
C231 a_n4866_1206# a_n7570_n1768# 0.255f
C232 a_n5100_n1638# a_n7570_n1768# 0.255f
C233 a_n5100_1206# a_n7570_n1768# 0.255f
C234 a_n5334_n1638# a_n7570_n1768# 0.255f
C235 a_n5334_1206# a_n7570_n1768# 0.255f
C236 a_n5568_n1638# a_n7570_n1768# 0.255f
C237 a_n5568_1206# a_n7570_n1768# 0.255f
C238 a_n5802_n1638# a_n7570_n1768# 0.255f
C239 a_n5802_1206# a_n7570_n1768# 0.255f
C240 a_n6036_n1638# a_n7570_n1768# 0.255f
C241 a_n6036_1206# a_n7570_n1768# 0.255f
C242 a_n6270_n1638# a_n7570_n1768# 0.255f
C243 a_n6270_1206# a_n7570_n1768# 0.255f
C244 a_n6504_n1638# a_n7570_n1768# 0.255f
C245 a_n6504_1206# a_n7570_n1768# 0.255f
C246 a_n6738_n1638# a_n7570_n1768# 0.255f
C247 a_n6738_1206# a_n7570_n1768# 0.255f
C248 a_n6972_n1638# a_n7570_n1768# 0.255f
C249 a_n6972_1206# a_n7570_n1768# 0.255f
C250 a_n7206_n1638# a_n7570_n1768# 0.255f
C251 a_n7206_1206# a_n7570_n1768# 0.255f
C252 a_n7440_n1638# a_n7570_n1768# 0.465f
C253 a_n7440_1206# a_n7570_n1768# 0.465f
.ends

.subckt IA_v4 VDD VSS G V1 V2 D0 D1 D2 D3 D4 D5 D6 D7 D8 D9 AVOUT1 AVOUT2 VOUT
Xx1 VDD x4/V2 D0 x1/m1_2124_1470# x1/m1_5470_410# x1/m1_2651_1472# x1/m1_3160_410#
+ x1/m1_4060_410# D3 D1 AVOUT1 D4 D2 G x1/m1_7940_410# RB_array_20
Xx3 VDD x6/V2 D5 x3/m1_2124_1470# x3/m1_5470_410# x3/m1_2651_1472# x3/m1_3160_410#
+ x3/m1_4060_410# D8 D6 VOUT D9 D7 G x3/m1_7940_410# RB_array_20
Xx2 VDD x5/V2 D0 x2/m1_2124_1470# x2/m1_5470_410# x2/m1_2651_1472# x2/m1_3160_410#
+ x2/m1_4060_410# D3 D1 AVOUT2 D4 D2 G x2/m1_7940_410# RB_array_20
Xx4 x4/V2 AVOUT1 x4/a_4864_8007# V2 x4/m1_4128_540# VDD x4/m1_5284_1188# x4/m1_4306_994#
+ x4/m3_5211_1261# VSS x4/m1_5053_7611# opamp
Xx5 x5/V2 AVOUT2 x5/a_4864_8007# V1 x5/m1_4128_540# VDD x5/m1_5284_1188# x5/m1_4306_994#
+ x5/m3_5211_1261# VSS x5/m1_5053_7611# opamp
Xx6 x6/V2 VOUT x6/a_4864_8007# x7/R1 x6/m1_4128_540# VDD x6/m1_5284_1188# x6/m1_4306_994#
+ x6/m3_5211_1261# VSS x6/m1_5053_7611# opamp
XXR1 x4/V2 x5/V2 x5/V2 x4/V2 x4/V2 x5/V2 x4/V2 x5/V2 x5/V2 x5/V2 x4/V2 x5/V2 x4/V2
+ x5/V2 x4/V2 x4/V2 x5/V2 x5/V2 x5/V2 x4/V2 x4/V2 x5/V2 x5/V2 x4/V2 x5/V2 x5/V2 x5/V2
+ x4/V2 x4/V2 x4/V2 x4/V2 x4/V2 x5/V2 x5/V2 x4/V2 x5/V2 x5/V2 x5/V2 x4/V2 x5/V2 x4/V2
+ x5/V2 x4/V2 x5/V2 x4/V2 x4/V2 x5/V2 x5/V2 x4/V2 x5/V2 x4/V2 x4/V2 x4/V2 x4/V2 x5/V2
+ x4/V2 x5/V2 x5/V2 x4/V2 x5/V2 x5/V2 x5/V2 x4/V2 x4/V2 x5/V2 x5/V2 x4/V2 x5/V2 x4/V2
+ x4/V2 x4/V2 x5/V2 x5/V2 x4/V2 x5/V2 x5/V2 x5/V2 x4/V2 x4/V2 x4/V2 x4/V2 x5/V2 x5/V2
+ x4/V2 x4/V2 x4/V2 x5/V2 x4/V2 x5/V2 x4/V2 x5/V2 x4/V2 x4/V2 x4/V2 x4/V2 x5/V2 x5/V2
+ x4/V2 x4/V2 x4/V2 x5/V2 x5/V2 x4/V2 x5/V2 G x5/V2 x5/V2 x5/V2 x4/V2 x5/V2 x4/V2
+ x4/V2 x5/V2 x5/V2 x4/V2 x4/V2 x4/V2 x5/V2 x5/V2 x4/V2 x5/V2 x5/V2 x4/V2 x4/V2 x5/V2
+ x5/V2 x4/V2 x4/V2 x5/V2 sky130_fd_pr__res_high_po_0p69_WX3C5M
Xx7 VDD x7/R1 D5 x7/m1_2124_1470# x7/m1_5470_410# x7/m1_2651_1472# x7/m1_3160_410#
+ x7/m1_4060_410# D8 D6 G D9 D7 G x7/m1_7940_410# RB_array_20
XXR2 x9/V2 x7/R1 x7/R1 x9/V2 x9/V2 x7/R1 x9/V2 x7/R1 x7/R1 x7/R1 x9/V2 x7/R1 x9/V2
+ x7/R1 x9/V2 x9/V2 x7/R1 x7/R1 x7/R1 x9/V2 x9/V2 x7/R1 x7/R1 x9/V2 x7/R1 x7/R1 x7/R1
+ x9/V2 x9/V2 x9/V2 x9/V2 x9/V2 x7/R1 x7/R1 x9/V2 x7/R1 x7/R1 x7/R1 x9/V2 x7/R1 x9/V2
+ x7/R1 x9/V2 x7/R1 x9/V2 x9/V2 x7/R1 x7/R1 x9/V2 x7/R1 x9/V2 x9/V2 x9/V2 x9/V2 x7/R1
+ x9/V2 x7/R1 x7/R1 x9/V2 x7/R1 x7/R1 x7/R1 x9/V2 x9/V2 x7/R1 x7/R1 x9/V2 x7/R1 x9/V2
+ x9/V2 x9/V2 x7/R1 x7/R1 x9/V2 x7/R1 x7/R1 x7/R1 x9/V2 x9/V2 x9/V2 x9/V2 x7/R1 x7/R1
+ x9/V2 x9/V2 x9/V2 x7/R1 x9/V2 x7/R1 x9/V2 x7/R1 x9/V2 x9/V2 x9/V2 x9/V2 x7/R1 x7/R1
+ x9/V2 x9/V2 x9/V2 x7/R1 x7/R1 x9/V2 x7/R1 G x7/R1 x7/R1 x7/R1 x9/V2 x7/R1 x9/V2
+ x9/V2 x7/R1 x7/R1 x9/V2 x9/V2 x9/V2 x7/R1 x7/R1 x9/V2 x7/R1 x7/R1 x9/V2 x9/V2 x7/R1
+ x7/R1 x9/V2 x9/V2 x7/R1 sky130_fd_pr__res_high_po_0p69_WX3C5M
Xx8 x8/V2 x8/V2 x8/a_4864_8007# AVOUT1 x8/m1_4128_540# VDD x8/m1_5284_1188# x8/m1_4306_994#
+ x8/m3_5211_1261# VSS x8/m1_5053_7611# opamp
Xx9 x9/V2 x9/V2 x9/a_4864_8007# AVOUT2 x9/m1_4128_540# VDD x9/m1_5284_1188# x9/m1_4306_994#
+ x9/m3_5211_1261# VSS x9/m1_5053_7611# opamp
XXR4 x8/V2 x6/V2 x6/V2 x8/V2 x8/V2 x6/V2 x8/V2 x6/V2 x6/V2 x6/V2 x8/V2 x6/V2 x8/V2
+ x6/V2 x8/V2 x8/V2 x6/V2 x6/V2 x6/V2 x8/V2 x8/V2 x6/V2 x6/V2 x8/V2 x6/V2 x6/V2 x6/V2
+ x8/V2 x8/V2 x8/V2 x8/V2 x8/V2 x6/V2 x6/V2 x8/V2 x6/V2 x6/V2 x6/V2 x8/V2 x6/V2 x8/V2
+ x6/V2 x8/V2 x6/V2 x8/V2 x8/V2 x6/V2 x6/V2 x8/V2 x6/V2 x8/V2 x8/V2 x8/V2 x8/V2 x6/V2
+ x8/V2 x6/V2 x6/V2 x8/V2 x6/V2 x6/V2 x6/V2 x8/V2 x8/V2 x6/V2 x6/V2 x8/V2 x6/V2 x8/V2
+ x8/V2 x8/V2 x6/V2 x6/V2 x8/V2 x6/V2 x6/V2 x6/V2 x8/V2 x8/V2 x8/V2 x8/V2 x6/V2 x6/V2
+ x8/V2 x8/V2 x8/V2 x6/V2 x8/V2 x6/V2 x8/V2 x6/V2 x8/V2 x8/V2 x8/V2 x8/V2 x6/V2 x6/V2
+ x8/V2 x8/V2 x8/V2 x6/V2 x6/V2 x8/V2 x6/V2 G x6/V2 x6/V2 x6/V2 x8/V2 x6/V2 x8/V2
+ x8/V2 x6/V2 x6/V2 x8/V2 x8/V2 x8/V2 x6/V2 x6/V2 x8/V2 x6/V2 x6/V2 x8/V2 x8/V2 x6/V2
+ x6/V2 x8/V2 x8/V2 x6/V2 sky130_fd_pr__res_high_po_0p69_WX3C5M
C0 x2/m1_7940_410# x7/m1_3160_410# 0.00253f
C1 AVOUT1 x5/V2 1.91f
C2 x4/V2 D1 0.0703f
C3 x4/m1_5284_1188# x5/m1_4128_540# 0.116f
C4 x8/m1_5053_7611# VDD 0.236f
C5 D0 D2 4.17e-25
C6 x3/m1_5470_410# D7 8.21e-20
C7 x5/m1_4306_994# AVOUT2 0.00888f
C8 x4/m1_4128_540# VDD 0.0784f
C9 x4/V2 D6 6.97e-20
C10 x6/V2 x6/a_4864_8007# 1.08f
C11 x2/m1_4060_410# D2 0.371f
C12 D0 D9 0.128f
C13 D5 VDD 0.302f
C14 x6/m1_5284_1188# VDD -0.00781f
C15 VDD x3/m1_3160_410# 1.98e-19
C16 x4/V2 x8/m1_5053_7611# 0.248f
C17 x6/m1_4128_540# x7/R1 0.0169f
C18 x4/V2 x4/m1_4128_540# 0.192f
C19 x2/m1_4060_410# D9 0.0424f
C20 x5/a_4864_8007# AVOUT1 0.0932f
C21 x4/V2 D5 8.21e-20
C22 x7/m1_5470_410# D9 0.113f
C23 D3 D2 0.00798f
C24 D5 x3/m1_2124_1470# 7.63e-19
C25 x9/m1_4128_540# x9/V2 0.0194f
C26 VOUT x9/V2 1.14f
C27 x9/a_4864_8007# x9/V2 0.162f
C28 D3 D9 0.126f
C29 x8/m3_5211_1261# AVOUT1 -0.0325f
C30 x9/m3_5211_1261# AVOUT2 -0.0333f
C31 x3/m1_2651_1472# VDD 2.09e-19
C32 V1 x5/V2 0.199f
C33 x6/V2 x9/V2 1.5f
C34 x8/m1_4306_994# AVOUT1 2.08f
C35 x3/m1_2651_1472# x3/m1_2124_1470# 3.55e-33
C36 VDD D4 3.74f
C37 x9/V2 x6/a_4864_8007# 0.136f
C38 x8/V2 x5/V2 3.14f
C39 x4/m3_5211_1261# VDD 0.00775f
C40 x5/a_4864_8007# V1 0.0336f
C41 x8/m1_5053_7611# x5/m1_5284_1188# 2.08e-20
C42 x5/m1_5053_7611# AVOUT1 0.0253f
C43 D2 D8 0.112f
C44 x4/V2 D4 0.071f
C45 D8 D9 5.8f
C46 x4/m3_5211_1261# x4/V2 0.0163f
C47 D4 x3/m1_2124_1470# 1.33e-19
C48 x5/m1_4306_994# x5/V2 0.122f
C49 D1 D2 0.244f
C50 x8/a_4864_8007# AVOUT1 -5.8e-19
C51 VOUT AVOUT1 0.0369f
C52 x9/m1_4128_540# AVOUT1 0.00295f
C53 D6 D2 0.112f
C54 D1 D9 0.128f
C55 x1/m1_5470_410# x1/m1_7940_410# -0.122f
C56 x1/m1_3160_410# AVOUT2 0.0165f
C57 x8/m1_5284_1188# AVOUT2 0.0242f
C58 D0 D7 0.112f
C59 x4/m1_5053_7611# VDD -0.236f
C60 x6/m1_4128_540# x9/m1_5053_7611# 0.251f
C61 D6 D9 0.128f
C62 x8/m3_5211_1261# x8/V2 0.00672f
C63 V2 VDD 0.133f
C64 x5/a_4864_8007# x5/m1_4306_994# -0.015f
C65 x6/m1_4128_540# VDD 0.118f
C66 x3/m1_5470_410# D8 0.00772f
C67 D5 D2 0.128f
C68 x7/m1_5470_410# D7 -3.46e-20
C69 x4/V2 x4/m1_5053_7611# 0.948f
C70 x8/m1_4128_540# AVOUT1 0.0796f
C71 x3/m1_7940_410# x7/R1 0.779f
C72 x5/m1_5053_7611# V1 0.00551f
C73 VOUT x9/m1_4306_994# 0.00253f
C74 D5 D9 0.129f
C75 x9/m1_4306_994# x9/a_4864_8007# -0.015f
C76 x4/V2 V2 0.199f
C77 x6/m1_4128_540# x4/V2 0.0527f
C78 D3 D7 0.108f
C79 x8/V2 x8/m1_4306_994# 0.0909f
C80 x3/m1_3160_410# D9 -0.00742f
C81 x7/R1 x5/V2 0.00553f
C82 VDD x7/m1_2651_1472# 5.3e-21
C83 x9/m1_5053_7611# AVOUT2 1.22f
C84 D0 x1/m1_2124_1470# -0.0315f
C85 x7/m1_2124_1470# D6 8.17e-20
C86 VDD AVOUT2 0.505f
C87 x8/V2 x8/a_4864_8007# 0.161f
C88 x2/m1_7940_410# x7/R1 0.0587f
C89 x8/V2 x9/m1_4128_540# 0.172f
C90 x4/a_4864_8007# VDD 0.0201f
C91 x7/m1_2124_1470# D5 0.0359f
C92 x4/V2 AVOUT2 0.34f
C93 x8/V2 x9/a_4864_8007# 0.384f
C94 x6/m1_5053_7611# VOUT -0.0477f
C95 D8 D7 5.38f
C96 D3 x2/m1_4060_410# -0.0252f
C97 x4/m1_5053_7611# x5/m1_4128_540# 0.251f
C98 D4 D9 0.148f
C99 x2/m1_2651_1472# x5/V2 2.84e-32
C100 x4/V2 x4/a_4864_8007# 1.16f
C101 x1/m1_3160_410# x5/V2 5.59e-19
C102 x8/V2 x6/V2 0.508f
C103 x1/m1_2651_1472# VDD 0.18f
C104 x6/m1_5053_7611# x6/V2 0.195f
C105 x8/V2 x8/m1_4128_540# 0.0193f
C106 D1 D7 0.111f
C107 x1/m1_7940_410# x6/V2 0.0587f
C108 x6/V2 x3/m1_4060_410# 0.34f
C109 x9/m1_4306_994# x9/V2 0.0905f
C110 x4/V2 x1/m1_2651_1472# 8.96e-20
C111 D6 D7 5.12f
C112 x6/m1_5053_7611# x6/a_4864_8007# -0.0112f
C113 D0 D8 0.112f
C114 D5 D7 0.112f
C115 x3/m1_3160_410# D7 -0.0172f
C116 x9/m3_5211_1261# VOUT 7.56e-19
C117 x7/m1_2124_1470# D4 1.33e-19
C118 x7/m1_5470_410# D8 0.327f
C119 AVOUT2 x5/m1_5284_1188# 0.0855f
C120 D0 D1 0.347f
C121 AVOUT2 x5/m1_4128_540# 0.00158f
C122 x6/m1_4306_994# VOUT 0.0139f
C123 D3 D8 0.108f
C124 D0 D6 0.112f
C125 x8/V2 x9/V2 0.00759f
C126 VDD x5/V2 5.66f
C127 x6/m1_5053_7611# x9/V2 2.57f
C128 VOUT x7/R1 1.42f
C129 x6/m1_4306_994# x6/V2 0.0347f
C130 D0 D5 0.127f
C131 x4/V2 x5/V2 0.7f
C132 x2/m1_7940_410# VDD 0.547f
C133 D9 x7/m1_2651_1472# 0.0126f
C134 D2 AVOUT2 0.611f
C135 x1/m1_5470_410# VDD 0.278f
C136 x6/V2 x7/R1 0.166f
C137 D3 D6 0.108f
C138 x5/a_4864_8007# VDD 0.0705f
C139 x2/m1_2651_1472# x2/m1_2124_1470# -0.0251f
C140 x6/m1_4306_994# x6/a_4864_8007# -2.59e-19
C141 D4 D7 0.115f
C142 x4/V2 x1/m1_5470_410# -0.00898f
C143 D3 D5 0.123f
C144 x4/V2 x5/a_4864_8007# 0.0335f
C145 x7/R1 x6/a_4864_8007# 0.189f
C146 x8/m1_5284_1188# x8/a_4864_8007# -0.00166f
C147 V1 AVOUT1 0.409f
C148 x8/m1_5284_1188# x9/m1_4128_540# 0.118f
C149 x8/m1_5284_1188# x9/a_4864_8007# 0.00572f
C150 V2 x4/m1_4306_994# -0.00251f
C151 x9/m3_5211_1261# x9/V2 0.00664f
C152 x8/m1_4306_994# VDD -0.00194f
C153 D1 D8 0.111f
C154 x2/m1_2651_1472# x2/m1_3160_410# -0.0129f
C155 x6/m1_4306_994# x9/V2 0.0128f
C156 x8/V2 AVOUT1 0.253f
C157 D6 D8 0.111f
C158 x5/m1_5284_1188# x5/V2 0.126f
C159 x5/V2 x5/m1_4128_540# 0.197f
C160 x5/m1_5053_7611# VDD -0.046f
C161 x2/m1_4060_410# D4 -0.00862f
C162 x7/R1 x9/V2 0.539f
C163 VDD x2/m1_5470_410# 0.291f
C164 x5/m1_4306_994# AVOUT1 0.0292f
C165 D5 D8 0.112f
C166 x2/m1_2124_1470# VDD 0.149f
C167 D6 D1 0.111f
C168 x3/m1_7940_410# D9 0.0078f
C169 x3/m1_3160_410# D8 -0.00742f
C170 x4/V2 x5/m1_5053_7611# 0.236f
C171 x8/V2 x9/m1_4306_994# 0.0139f
C172 D3 D4 -0.00199f
C173 x9/m1_5053_7611# VOUT 0.00204f
C174 x5/a_4864_8007# x5/m1_5284_1188# -0.00166f
C175 x9/m1_5053_7611# x9/m1_4128_540# -0.00132f
C176 VDD x8/a_4864_8007# 0.112f
C177 x9/m1_5053_7611# x9/a_4864_8007# -0.00138f
C178 x5/a_4864_8007# x5/m1_4128_540# -0.00634f
C179 VDD x9/m1_4128_540# 0.201f
C180 VOUT VDD 0.0955f
C181 D5 D1 0.127f
C182 x1/m1_4060_410# VDD 0.224f
C183 VDD x9/a_4864_8007# 0.112f
C184 D2 x5/V2 0.197f
C185 x4/a_4864_8007# x4/m1_4306_994# -0.015f
C186 x4/V2 x8/a_4864_8007# 0.0335f
C187 x9/m1_5053_7611# x6/V2 0.033f
C188 D7 x7/m1_2651_1472# 2.24e-20
C189 D6 D5 4.98f
C190 x5/m3_5211_1261# AVOUT2 0.00626f
C191 D9 x5/V2 0.123f
C192 x4/V2 x9/m1_4128_540# 0.0515f
C193 VDD x6/V2 4.94f
C194 D6 x3/m1_3160_410# 0.00749f
C195 x8/m1_5284_1188# x9/V2 0.0252f
C196 x4/V2 x9/a_4864_8007# 0.0335f
C197 x4/V2 x1/m1_4060_410# -0.00329f
C198 x8/m1_4128_540# VDD 0.224f
C199 x2/m1_3160_410# VDD 0.196f
C200 x1/m1_5470_410# D2 7.1e-20
C201 x9/m1_5053_7611# x6/a_4864_8007# 0.0605f
C202 x4/V2 x6/V2 0.551f
C203 x8/m1_4306_994# x5/m1_5284_1188# 0.129f
C204 D5 x3/m1_3160_410# 4.76e-19
C205 x5/m1_4306_994# V1 -0.00251f
C206 x2/m1_7940_410# D9 0.188f
C207 VDD x6/a_4864_8007# -0.017f
C208 x4/m1_5053_7611# x4/m1_5284_1188# -0.00274f
C209 x4/V2 x8/m1_4128_540# 0.0532f
C210 x6/V2 x3/m1_2124_1470# 5.38e-19
C211 D4 D8 0.115f
C212 x3/m1_2651_1472# D6 4.73e-19
C213 x4/V2 x6/a_4864_8007# 0.0305f
C214 x5/m1_5053_7611# x5/m1_4128_540# -0.00124f
C215 x6/m1_4128_540# x9/m1_5284_1188# 0.116f
C216 x3/m1_2651_1472# D5 0.0354f
C217 D0 AVOUT2 0.525f
C218 D6 D4 0.115f
C219 x9/m1_5053_7611# x9/V2 0.39f
C220 x8/a_4864_8007# x5/m1_5284_1188# 0.00572f
C221 VDD x9/V2 2.98f
C222 x1/m1_2124_1470# AVOUT2 0.00826f
C223 x2/m1_7940_410# x7/m1_2124_1470# 0.0514f
C224 D5 D4 0.133f
C225 x8/m1_5284_1188# AVOUT1 0.0237f
C226 D3 AVOUT2 0.705f
C227 x4/V2 x9/V2 0.112f
C228 D0 x1/m1_2651_1472# 0.00477f
C229 AVOUT2 x4/m1_5284_1188# 3.25e-20
C230 x8/V2 x9/m3_5211_1261# 5.32e-20
C231 x8/m1_4128_540# x5/m1_5284_1188# 0.118f
C232 x5/m3_5211_1261# x5/V2 0.0161f
C233 x2/m1_5470_410# D9 0.0828f
C234 x2/m1_2124_1470# D9 0.0126f
C235 x9/m1_5284_1188# AVOUT2 7.6e-20
C236 x4/a_4864_8007# x4/m1_5284_1188# -0.00166f
C237 D7 x5/V2 0.104f
C238 x1/m1_4060_410# D2 -9.41e-19
C239 x8/m1_5284_1188# x9/m1_4306_994# 0.129f
C240 x3/m1_2651_1472# D4 5.48e-20
C241 x4/m1_5053_7611# x4/m1_4128_540# -0.00195f
C242 x6/m1_5053_7611# x7/R1 0.771f
C243 V2 x4/m1_4128_540# 0.00448f
C244 x2/m1_7940_410# D7 0.0346f
C245 x2/m1_3160_410# D2 0.0412f
C246 x6/V2 D9 0.123f
C247 x2/m1_3160_410# D9 0.0228f
C248 VDD AVOUT1 0.313f
C249 D0 x5/V2 -3.64e-19
C250 D6 x7/m1_2651_1472# 0.0168f
C251 D1 AVOUT2 0.553f
C252 x4/V2 AVOUT1 0.295f
C253 x2/m1_4060_410# x5/V2 0.613f
C254 x8/V2 x8/m1_5284_1188# 0.344f
C255 x9/m1_5053_7611# x9/m1_4306_994# -0.626f
C256 x3/m1_5470_410# x6/V2 2.58e-20
C257 D5 x7/m1_2651_1472# 0.423f
C258 VDD x9/m1_4306_994# -0.00194f
C259 x8/m1_5053_7611# AVOUT2 0.0247f
C260 D3 x5/V2 1.15f
C261 x4/m1_5284_1188# x5/V2 0.0389f
C262 D5 AVOUT2 0.55f
C263 D1 x1/m1_2651_1472# -0.0116f
C264 x6/m1_4306_994# x7/R1 0.00314f
C265 x4/a_4864_8007# x4/m1_4128_540# -0.0213f
C266 VDD V1 1.99f
C267 D3 x1/m1_5470_410# -0.0126f
C268 x5/a_4864_8007# x4/m1_5284_1188# 0.00551f
C269 x4/V2 V1 0.27f
C270 x8/V2 x9/m1_5053_7611# 0.662f
C271 x6/m1_5053_7611# x9/m1_5053_7611# 0.181f
C272 x5/m1_5284_1188# AVOUT1 0.0238f
C273 x8/V2 VDD 1.52f
C274 AVOUT1 x5/m1_4128_540# 0.204f
C275 x6/m1_5053_7611# VDD -0.276f
C276 x7/m1_4060_410# D9 0.0424f
C277 D8 x5/V2 0.104f
C278 D4 x7/m1_2651_1472# 5.48e-20
C279 x1/m1_7940_410# VDD 0.519f
C280 x6/V2 D7 0.165f
C281 x4/V2 x8/V2 0.783f
C282 x4/V2 x6/m1_5053_7611# 0.16f
C283 AVOUT2 D4 1.11f
C284 x5/m1_4306_994# VDD -0.00155f
C285 D0 x2/m1_2124_1470# 0.037f
C286 x7/m1_3160_410# D9 0.0228f
C287 D1 x5/V2 6.38e-22
C288 x4/V2 x1/m1_7940_410# -0.00872f
C289 x2/m1_4060_410# x2/m1_5470_410# -0.098f
C290 x2/m1_7940_410# D8 0.0346f
C291 x1/m1_7940_410# x3/m1_2124_1470# 0.0514f
C292 D6 x5/V2 0.104f
C293 x4/m3_5211_1261# x4/a_4864_8007# -0.00142f
C294 x8/m1_5053_7611# x5/V2 4.5e-19
C295 x5/m1_5053_7611# x4/m1_5284_1188# 2.08e-20
C296 D3 x2/m1_5470_410# 0.293f
C297 D5 x5/V2 0.119f
C298 V1 x5/m1_4128_540# 0.0262f
C299 x2/m1_7940_410# D6 0.0346f
C300 D0 x2/m1_3160_410# 6.29e-19
C301 D3 x1/m1_4060_410# -0.0278f
C302 x6/m1_4306_994# VDD 0.00401f
C303 x2/m1_3160_410# x2/m1_4060_410# -0.00924f
C304 x2/m1_7940_410# D5 0.0379f
C305 x7/m1_7940_410# x7/R1 0.99f
C306 x4/m1_5053_7611# x4/a_4864_8007# -0.00354f
C307 x8/V2 x5/m1_5284_1188# 0.0252f
C308 VOUT x6/m3_5211_1261# 0.0102f
C309 x9/m1_5284_1188# VOUT 0.0226f
C310 x9/m1_5284_1188# x9/a_4864_8007# -0.00166f
C311 x4/a_4864_8007# V2 0.00147f
C312 VDD x7/R1 1.63f
C313 x6/V2 x6/m3_5211_1261# 0.0101f
C314 x9/m1_5284_1188# x6/V2 0.054f
C315 x7/m1_4060_410# D7 0.368f
C316 x8/m1_4306_994# x8/m1_5053_7611# -0.627f
C317 D4 x5/V2 0.178f
C318 x6/a_4864_8007# x6/m3_5211_1261# -0.00131f
C319 x9/m1_5284_1188# x6/a_4864_8007# 0.00551f
C320 x4/m1_4306_994# AVOUT1 0.0138f
C321 x2/m1_2651_1472# VDD 0.164f
C322 x9/m1_5053_7611# x8/m1_5284_1188# 2.08e-20
C323 x7/m1_3160_410# D7 0.0234f
C324 x8/m1_5053_7611# x5/m1_5053_7611# 0.198f
C325 x1/m1_3160_410# VDD 0.206f
C326 x8/m1_5284_1188# VDD -0.0958f
C327 x6/V2 D8 0.102f
C328 x2/m1_7940_410# D4 0.448f
C329 x1/m1_7940_410# D9 0.0346f
C330 x5/m3_5211_1261# AVOUT1 0.0068f
C331 D9 x3/m1_4060_410# -0.0064f
C332 x1/m1_5470_410# D4 -0.0325f
C333 x1/m1_4060_410# D1 2.24e-19
C334 x4/V2 x1/m1_3160_410# 4.41e-20
C335 x8/m1_5053_7611# x8/a_4864_8007# -0.00138f
C336 x8/m1_5053_7611# x9/m1_4128_540# 0.251f
C337 x1/m1_2651_1472# AVOUT2 0.00829f
C338 x8/m1_5053_7611# x9/a_4864_8007# 0.0618f
C339 x9/V2 x6/m3_5211_1261# 5.32e-20
C340 x9/m1_5284_1188# x9/V2 0.341f
C341 x2/m1_3160_410# D1 0.42f
C342 D6 x6/V2 0.0361f
C343 x6/m1_5284_1188# VOUT 0.15f
C344 x4/m1_4306_994# V1 0.00225f
C345 x8/m1_5053_7611# x8/m1_4128_540# -0.00132f
C346 D5 x6/V2 0.063f
C347 x5/a_4864_8007# x4/m1_5053_7611# 0.0587f
C348 x9/m1_5053_7611# VDD 0.0851f
C349 x3/m1_3160_410# x6/V2 0.557f
C350 x4/V2 x9/m1_5053_7611# 0.239f
C351 x2/m1_5470_410# D4 0.041f
C352 x6/m1_5284_1188# x6/a_4864_8007# -5.52e-19
C353 x4/V2 VDD 8.38f
C354 x7/R1 D9 0.137f
C355 VDD x3/m1_2124_1470# 7.88e-19
C356 x3/m1_2651_1472# x6/V2 -0.00694f
C357 AVOUT2 x5/V2 0.557f
C358 x4/m1_5284_1188# AVOUT1 0.103f
C359 x2/m1_7940_410# x7/m1_2651_1472# 1.19e-19
C360 x1/m1_4060_410# D4 -0.00862f
C361 x7/m1_4060_410# D8 0.0291f
C362 x1/m1_7940_410# D7 0.0346f
C363 D7 x3/m1_4060_410# 0.00157f
C364 x2/m1_2651_1472# D2 9.01e-22
C365 x1/m1_5470_410# AVOUT2 0.742f
C366 x4/m1_5053_7611# x5/m1_5053_7611# 0.197f
C367 D4 x6/V2 8.91e-19
C368 x5/a_4864_8007# AVOUT2 -0.00792f
C369 x1/m1_3160_410# D2 -0.00573f
C370 x6/m1_5284_1188# x9/V2 0.00765f
C371 x2/m1_2651_1472# D9 0.0126f
C372 D6 x7/m1_4060_410# 1.64e-19
C373 x8/m3_5211_1261# AVOUT2 0.00644f
C374 VDD x5/m1_5284_1188# -0.0331f
C375 VDD x5/m1_4128_540# 0.197f
C376 D5 x7/m1_4060_410# -7.28e-21
C377 V1 x4/m1_5284_1188# 0.0196f
C378 x7/m1_3160_410# D6 0.394f
C379 x6/m1_4128_540# VOUT 0.0402f
C380 x8/m1_4306_994# AVOUT2 0.0551f
C381 x4/V2 x5/m1_4128_540# 0.0538f
C382 x6/m1_4128_540# x6/V2 0.203f
C383 x7/m1_3160_410# D5 0.00102f
C384 x5/m1_5053_7611# AVOUT2 -0.0011f
C385 x8/m1_5053_7611# AVOUT1 1.25f
C386 D3 x1/m1_7940_410# -1.11e-20
C387 D2 VDD 1.46f
C388 x7/m1_7940_410# D9 0.462f
C389 x4/m1_4128_540# AVOUT1 0.0348f
C390 x6/m1_4128_540# x6/a_4864_8007# -0.00333f
C391 x7/R1 D7 0.0157f
C392 VDD D9 0.254f
C393 x6/m1_5053_7611# x9/m1_5284_1188# 2.08e-20
C394 x4/V2 D2 0.0705f
C395 x5/m1_4306_994# x4/m1_5284_1188# 0.129f
C396 x8/a_4864_8007# AVOUT2 0.462f
C397 x9/m1_4128_540# AVOUT2 0.116f
C398 VOUT AVOUT2 0.0201f
C399 x2/m1_7940_410# x5/V2 -1.13e-31
C400 x1/m1_4060_410# AVOUT2 0.022f
C401 AVOUT2 x9/a_4864_8007# 7.79e-19
C402 x1/m1_5470_410# x5/V2 0.349f
C403 x5/a_4864_8007# x5/V2 1.16f
C404 x8/m1_4128_540# AVOUT2 0.25f
C405 x6/m1_4128_540# x9/V2 0.205f
C406 x1/m1_7940_410# D8 0.0346f
C407 D8 x3/m1_4060_410# -0.0058f
C408 x4/m1_4128_540# V1 0.136f
C409 x7/m1_2124_1470# VDD 0.00904f
C410 x4/m3_5211_1261# AVOUT1 0.00702f
C411 x9/m1_5284_1188# x6/m1_4306_994# 0.129f
C412 x8/V2 x8/m1_5053_7611# 0.391f
C413 D6 x3/m1_4060_410# 2.24e-19
C414 D6 x1/m1_7940_410# 0.0346f
C415 x4/m1_4306_994# VDD 0.0222f
C416 x5/m1_5053_7611# x5/V2 0.741f
C417 D0 x2/m1_2651_1472# 0.489f
C418 x7/R1 x6/m3_5211_1261# 3.23e-19
C419 D0 x1/m1_3160_410# 4.76e-19
C420 x2/m1_5470_410# x5/V2 0.254f
C421 x9/m1_5284_1188# x7/R1 7.44e-20
C422 x6/m1_5053_7611# x6/m1_5284_1188# -0.00236f
C423 D5 x1/m1_7940_410# 0.0355f
C424 x4/V2 x4/m1_4306_994# 0.123f
C425 AVOUT2 x9/V2 0.219f
C426 x1/m1_7940_410# x3/m1_3160_410# 0.00253f
C427 x3/m1_3160_410# x3/m1_4060_410# -0.116f
C428 VDD D7 0.193f
C429 x5/a_4864_8007# x5/m1_5053_7611# -0.00316f
C430 x4/m1_5053_7611# AVOUT1 -0.0659f
C431 x1/m1_4060_410# x5/V2 0.67f
C432 V2 AVOUT1 0.00262f
C433 D2 D9 0.13f
C434 x4/V2 D7 6.97e-20
C435 x4/m3_5211_1261# V1 2.71e-19
C436 x7/R1 D8 0.0218f
C437 x6/V2 x5/V2 0.508f
C438 x3/m1_2651_1472# x1/m1_7940_410# 1.19e-19
C439 x8/m1_4128_540# x5/V2 5.49e-19
C440 x2/m1_3160_410# x5/V2 1.37e-20
C441 x1/m1_5470_410# x1/m1_4060_410# -0.121f
C442 D0 VDD 1.25f
C443 D6 x7/R1 0.0104f
C444 x1/m1_7940_410# D4 -0.0234f
C445 x2/m1_4060_410# VDD 0.218f
C446 x4/m1_5053_7611# V1 0.747f
C447 VDD x1/m1_2124_1470# 0.151f
C448 x3/m1_5470_410# D9 6.59e-19
C449 D0 x4/V2 0.0701f
C450 AVOUT2 AVOUT1 1.09f
C451 x8/m1_4306_994# x8/a_4864_8007# -0.015f
C452 D5 x7/R1 -4.54e-20
C453 V2 V1 0.0641f
C454 x6/m1_5284_1188# x7/R1 0.0337f
C455 D3 VDD 2.3f
C456 x4/V2 x1/m1_2124_1470# 0.0518f
C457 x2/m1_2651_1472# D1 0.0265f
C458 x4/a_4864_8007# AVOUT1 -0.00756f
C459 VDD x4/m1_5284_1188# -0.0358f
C460 x7/m1_2124_1470# D9 0.0126f
C461 x1/m1_3160_410# D1 0.00239f
C462 x9/m1_5053_7611# x9/m1_5284_1188# -0.00704f
C463 x5/m1_5053_7611# x8/a_4864_8007# 0.0618f
C464 D3 x4/V2 0.0711f
C465 x9/m1_5284_1188# VDD -0.0958f
C466 x9/m1_4306_994# AVOUT2 2.15f
C467 x4/V2 x4/m1_5284_1188# 0.129f
C468 x6/m1_4128_540# x6/m1_5053_7611# -0.00104f
C469 x8/m1_5053_7611# x8/m1_5284_1188# -0.00704f
C470 x8/m1_4128_540# x5/m1_5053_7611# 0.257f
C471 x7/m1_7940_410# D8 -1.6e-19
C472 VOUT x9/m1_4128_540# 0.00868f
C473 AVOUT2 V1 -2.31e-19
C474 x9/m1_4128_540# x9/a_4864_8007# -0.00709f
C475 D2 D7 0.112f
C476 VDD D8 0.191f
C477 D4 x7/R1 8.91e-19
C478 D7 D9 0.129f
C479 x4/a_4864_8007# V1 0.548f
C480 VOUT x6/V2 0.601f
C481 x8/m1_4128_540# x8/a_4864_8007# -0.0068f
C482 x4/V2 D8 6.97e-20
C483 x8/V2 AVOUT2 0.619f
C484 D1 VDD 1.12f
C485 x1/m1_7940_410# AVOUT2 0.583f
C486 D6 VDD 0.199f
C487 x8/m1_5053_7611# x9/m1_5053_7611# 0.184f
C488 dw_n60_n20# VSS 0.339p **FLOATING
C489 x8/V2 VSS 30.1f
C490 x9/m3_5211_1261# VSS 0.916f
C491 x9/m1_5053_7611# VSS 4.5f
C492 x9/m1_5284_1188# VSS 4.46f
C493 x9/m1_4306_994# VSS 5.89f
C494 x9/a_4864_8007# VSS 5.11f
C495 x9/m1_4128_540# VSS 2.64f
C496 x8/m3_5211_1261# VSS 0.907f
C497 x8/m1_5053_7611# VSS 4.51f
C498 x8/m1_5284_1188# VSS 4.48f
C499 x8/m1_4306_994# VSS 5.86f
C500 x8/a_4864_8007# VSS 5.07f
C501 x8/m1_4128_540# VSS 2.6f
C502 x9/V2 VSS 27.9f
C503 x7/R1 VSS 36.8f
C504 x7/m1_7940_410# VSS 6.21f
C505 D9 VSS 26.1f
C506 D7 VSS 11.3f
C507 D8 VSS 16.6f
C508 D6 VSS 8.14f
C509 D5 VSS 7.8f
C510 x7/m1_4060_410# VSS 2.26f
C511 x7/m1_5470_410# VSS 3.44f
C512 x7/m1_3160_410# VSS 1.68f
C513 x7/m1_2124_1470# VSS 1.08f
C514 x7/m1_2651_1472# VSS 1f
C515 x6/m3_5211_1261# VSS 0.892f
C516 x6/m1_5053_7611# VSS 4.53f
C517 x6/m1_5284_1188# VSS 4.44f
C518 x6/m1_4306_994# VSS 5.85f
C519 x6/a_4864_8007# VSS 4.81f
C520 x6/m1_4128_540# VSS 2.57f
C521 x5/m3_5211_1261# VSS 0.884f
C522 x5/m1_5053_7611# VSS 4.5f
C523 x5/m1_5284_1188# VSS 4.46f
C524 V1 VSS 1.04f
C525 x5/m1_4306_994# VSS 5.81f
C526 x5/a_4864_8007# VSS 4.8f
C527 x5/m1_4128_540# VSS 2.53f
C528 x4/m3_5211_1261# VSS 0.88f
C529 VDD VSS 0.228p
C530 x4/m1_5053_7611# VSS 4.56f
C531 x4/m1_5284_1188# VSS 4.43f
C532 V2 VSS 1.01f
C533 x4/m1_4306_994# VSS 5.78f
C534 x4/a_4864_8007# VSS 4.83f
C535 x4/m1_4128_540# VSS 2.51f
C536 x5/V2 VSS 41.8f
C537 x2/m1_7940_410# VSS 6.21f
C538 D4 VSS 17.8f
C539 D2 VSS 5.9f
C540 D3 VSS 10.4f
C541 D1 VSS 3.57f
C542 D0 VSS 2.7f
C543 x2/m1_4060_410# VSS 2.12f
C544 x2/m1_5470_410# VSS 3.36f
C545 x2/m1_3160_410# VSS 1.66f
C546 AVOUT2 VSS 20.5f
C547 x2/m1_2124_1470# VSS 1.08f
C548 x2/m1_2651_1472# VSS 0.966f
C549 x6/V2 VSS 39.4f
C550 x3/m1_7940_410# VSS 6.27f
C551 x3/m1_4060_410# VSS 2.22f
C552 x3/m1_5470_410# VSS 3.48f
C553 x3/m1_3160_410# VSS 1.59f
C554 VOUT VSS 18.7f
C555 x3/m1_2124_1470# VSS 1.11f
C556 x3/m1_2651_1472# VSS 1.01f
C557 x4/V2 VSS 35.8f
C558 x1/m1_7940_410# VSS 6.21f
C559 x1/m1_4060_410# VSS 2.12f
C560 x1/m1_5470_410# VSS 3.22f
C561 x1/m1_3160_410# VSS 1.69f
C562 AVOUT1 VSS 17.5f
C563 x1/m1_2124_1470# VSS 1.09f
C564 x1/m1_2651_1472# VSS 1f
.ends

