* SPICE3 file created from RB_array_20.ext - technology: sky130A

.subckt sky130_fd_pr__res_high_po_0p69_JKKHRG a_n199_n1768# a_n69_1206# a_n69_n1638#
X0 a_n69_1206# a_n69_n1638# a_n199_n1768# sky130_fd_pr__res_high_po_0p69 l=12.1
C0 a_n69_n1638# a_n199_n1768# 0.675f
C1 a_n69_1206# a_n199_n1768# 0.675f
.ends

.subckt sky130_fd_pr__res_high_po_0p69_Z3RMRJ a_48_1206# a_n186_n1638# a_n186_1206#
+ a_n316_n1768# a_48_n1638#
X0 a_48_1206# a_48_n1638# a_n316_n1768# sky130_fd_pr__res_high_po_0p69 l=12.1
X1 a_n186_1206# a_n186_n1638# a_n316_n1768# sky130_fd_pr__res_high_po_0p69 l=12.1
C0 a_48_1206# a_n186_1206# 0.296f
C1 a_n186_n1638# a_48_n1638# 0.296f
C2 a_48_n1638# a_n316_n1768# 0.465f
C3 a_48_1206# a_n316_n1768# 0.465f
C4 a_n186_n1638# a_n316_n1768# 0.465f
C5 a_n186_1206# a_n316_n1768# 0.465f
.ends

.subckt sky130_fd_pr__res_high_po_0p69_Z3RMR6 a_516_n1638# a_48_1206# a_n654_1206#
+ a_n888_1206# a_n186_n1638# a_n186_1206# a_750_1206# a_n654_n1638# a_282_1206# a_282_n1638#
+ a_48_n1638# a_750_n1638# a_n420_n1638# a_516_1206# a_n1018_n1768# a_n420_1206# a_n888_n1638#
X0 a_n420_1206# a_n420_n1638# a_n1018_n1768# sky130_fd_pr__res_high_po_0p69 l=12.1
X1 a_48_1206# a_48_n1638# a_n1018_n1768# sky130_fd_pr__res_high_po_0p69 l=12.1
X2 a_750_1206# a_750_n1638# a_n1018_n1768# sky130_fd_pr__res_high_po_0p69 l=12.1
X3 a_n888_1206# a_n888_n1638# a_n1018_n1768# sky130_fd_pr__res_high_po_0p69 l=12.1
X4 a_282_1206# a_282_n1638# a_n1018_n1768# sky130_fd_pr__res_high_po_0p69 l=12.1
X5 a_n654_1206# a_n654_n1638# a_n1018_n1768# sky130_fd_pr__res_high_po_0p69 l=12.1
X6 a_n186_1206# a_n186_n1638# a_n1018_n1768# sky130_fd_pr__res_high_po_0p69 l=12.1
X7 a_516_1206# a_516_n1638# a_n1018_n1768# sky130_fd_pr__res_high_po_0p69 l=12.1
C0 a_48_n1638# a_n186_n1638# 0.296f
C1 a_n186_1206# a_n420_1206# 0.296f
C2 a_750_n1638# a_516_n1638# 0.296f
C3 a_n420_n1638# a_n654_n1638# 0.296f
C4 a_282_1206# a_516_1206# 0.296f
C5 a_48_n1638# a_282_n1638# 0.296f
C6 a_750_1206# a_516_1206# 0.296f
C7 a_516_n1638# a_282_n1638# 0.296f
C8 a_n654_1206# a_n888_1206# 0.296f
C9 a_n654_1206# a_n420_1206# 0.296f
C10 a_n888_n1638# a_n654_n1638# 0.296f
C11 a_48_1206# a_n186_1206# 0.296f
C12 a_282_1206# a_48_1206# 0.296f
C13 a_n186_n1638# a_n420_n1638# 0.296f
C14 a_750_n1638# a_n1018_n1768# 0.465f
C15 a_750_1206# a_n1018_n1768# 0.465f
C16 a_516_n1638# a_n1018_n1768# 0.255f
C17 a_516_1206# a_n1018_n1768# 0.255f
C18 a_282_n1638# a_n1018_n1768# 0.255f
C19 a_282_1206# a_n1018_n1768# 0.255f
C20 a_48_n1638# a_n1018_n1768# 0.255f
C21 a_48_1206# a_n1018_n1768# 0.255f
C22 a_n186_n1638# a_n1018_n1768# 0.255f
C23 a_n186_1206# a_n1018_n1768# 0.255f
C24 a_n420_n1638# a_n1018_n1768# 0.255f
C25 a_n420_1206# a_n1018_n1768# 0.255f
C26 a_n654_n1638# a_n1018_n1768# 0.255f
C27 a_n654_1206# a_n1018_n1768# 0.255f
C28 a_n888_n1638# a_n1018_n1768# 0.465f
C29 a_n888_1206# a_n1018_n1768# 0.465f
.ends

.subckt sky130_fd_pr__res_high_po_0p69_YMHKRJ a_48_1206# a_n550_n1768# a_n186_n1638#
+ a_n186_1206# a_282_1206# a_282_n1638# a_48_n1638# a_n420_n1638# a_n420_1206#
X0 a_n420_1206# a_n420_n1638# a_n550_n1768# sky130_fd_pr__res_high_po_0p69 l=12.1
X1 a_48_1206# a_48_n1638# a_n550_n1768# sky130_fd_pr__res_high_po_0p69 l=12.1
X2 a_282_1206# a_282_n1638# a_n550_n1768# sky130_fd_pr__res_high_po_0p69 l=12.1
X3 a_n186_1206# a_n186_n1638# a_n550_n1768# sky130_fd_pr__res_high_po_0p69 l=12.1
C0 a_n186_n1638# a_n420_n1638# 0.296f
C1 a_n186_n1638# a_48_n1638# 0.296f
C2 a_n186_1206# a_n420_1206# 0.296f
C3 a_n186_1206# a_48_1206# 0.296f
C4 a_282_n1638# a_48_n1638# 0.296f
C5 a_282_1206# a_48_1206# 0.296f
C6 a_282_n1638# a_n550_n1768# 0.465f
C7 a_282_1206# a_n550_n1768# 0.465f
C8 a_48_n1638# a_n550_n1768# 0.255f
C9 a_48_1206# a_n550_n1768# 0.255f
C10 a_n186_n1638# a_n550_n1768# 0.255f
C11 a_n186_1206# a_n550_n1768# 0.255f
C12 a_n420_n1638# a_n550_n1768# 0.465f
C13 a_n420_1206# a_n550_n1768# 0.465f
.ends

.subckt sky130_fd_pr__res_high_po_0p69_HBQF5Z a_516_n1638# a_48_1206# a_n654_1206#
+ a_n888_1206# a_1452_1206# a_n1122_n1638# a_1452_n1638# a_n186_n1638# a_n186_1206#
+ a_n1954_n1768# a_1686_1206# a_750_1206# a_n654_n1638# a_n1590_1206# a_984_n1638#
+ a_984_1206# a_n1824_1206# a_n1590_n1638# a_1218_n1638# a_282_1206# a_n1122_1206#
+ a_1218_1206# a_282_n1638# a_48_n1638# a_750_n1638# a_n420_n1638# a_n1356_1206# a_516_1206#
+ a_n1356_n1638# a_1686_n1638# a_n420_1206# a_n1824_n1638# a_n888_n1638#
X0 a_n420_1206# a_n420_n1638# a_n1954_n1768# sky130_fd_pr__res_high_po_0p69 l=12.1
X1 a_1452_1206# a_1452_n1638# a_n1954_n1768# sky130_fd_pr__res_high_po_0p69 l=12.1
X2 a_n1824_1206# a_n1824_n1638# a_n1954_n1768# sky130_fd_pr__res_high_po_0p69 l=12.1
X3 a_n1590_1206# a_n1590_n1638# a_n1954_n1768# sky130_fd_pr__res_high_po_0p69 l=12.1
X4 a_48_1206# a_48_n1638# a_n1954_n1768# sky130_fd_pr__res_high_po_0p69 l=12.1
X5 a_984_1206# a_984_n1638# a_n1954_n1768# sky130_fd_pr__res_high_po_0p69 l=12.1
X6 a_n1356_1206# a_n1356_n1638# a_n1954_n1768# sky130_fd_pr__res_high_po_0p69 l=12.1
X7 a_1218_1206# a_1218_n1638# a_n1954_n1768# sky130_fd_pr__res_high_po_0p69 l=12.1
X8 a_750_1206# a_750_n1638# a_n1954_n1768# sky130_fd_pr__res_high_po_0p69 l=12.1
X9 a_n1122_1206# a_n1122_n1638# a_n1954_n1768# sky130_fd_pr__res_high_po_0p69 l=12.1
X10 a_n888_1206# a_n888_n1638# a_n1954_n1768# sky130_fd_pr__res_high_po_0p69 l=12.1
X11 a_282_1206# a_282_n1638# a_n1954_n1768# sky130_fd_pr__res_high_po_0p69 l=12.1
X12 a_n654_1206# a_n654_n1638# a_n1954_n1768# sky130_fd_pr__res_high_po_0p69 l=12.1
X13 a_n186_1206# a_n186_n1638# a_n1954_n1768# sky130_fd_pr__res_high_po_0p69 l=12.1
X14 a_516_1206# a_516_n1638# a_n1954_n1768# sky130_fd_pr__res_high_po_0p69 l=12.1
X15 a_1686_1206# a_1686_n1638# a_n1954_n1768# sky130_fd_pr__res_high_po_0p69 l=12.1
C0 a_n420_1206# a_n186_1206# 0.296f
C1 a_n654_n1638# a_n420_n1638# 0.296f
C2 a_516_1206# a_282_1206# 0.296f
C3 a_n888_1206# a_n654_1206# 0.296f
C4 a_282_n1638# a_48_n1638# 0.296f
C5 a_n1122_n1638# a_n888_n1638# 0.296f
C6 a_n420_1206# a_n654_1206# 0.296f
C7 a_1686_n1638# a_1452_n1638# 0.296f
C8 a_n654_n1638# a_n888_n1638# 0.296f
C9 a_48_1206# a_282_1206# 0.296f
C10 a_n186_n1638# a_48_n1638# 0.296f
C11 a_n1590_n1638# a_n1356_n1638# 0.296f
C12 a_48_1206# a_n186_1206# 0.296f
C13 a_n186_n1638# a_n420_n1638# 0.296f
C14 a_n1356_1206# a_n1590_1206# 0.296f
C15 a_1218_1206# a_984_1206# 0.296f
C16 a_984_n1638# a_750_n1638# 0.296f
C17 a_750_1206# a_516_1206# 0.296f
C18 a_1452_1206# a_1686_1206# 0.296f
C19 a_516_n1638# a_282_n1638# 0.296f
C20 a_1218_n1638# a_1452_n1638# 0.296f
C21 a_1452_1206# a_1218_1206# 0.296f
C22 a_750_1206# a_984_1206# 0.296f
C23 a_1218_n1638# a_984_n1638# 0.296f
C24 a_n888_1206# a_n1122_1206# 0.296f
C25 a_516_n1638# a_750_n1638# 0.296f
C26 a_n1590_n1638# a_n1824_n1638# 0.296f
C27 a_n1122_n1638# a_n1356_n1638# 0.296f
C28 a_n1356_1206# a_n1122_1206# 0.296f
C29 a_n1590_1206# a_n1824_1206# 0.296f
C30 a_1686_n1638# a_n1954_n1768# 0.465f
C31 a_1686_1206# a_n1954_n1768# 0.465f
C32 a_1452_n1638# a_n1954_n1768# 0.255f
C33 a_1452_1206# a_n1954_n1768# 0.255f
C34 a_1218_n1638# a_n1954_n1768# 0.255f
C35 a_1218_1206# a_n1954_n1768# 0.255f
C36 a_984_n1638# a_n1954_n1768# 0.255f
C37 a_984_1206# a_n1954_n1768# 0.255f
C38 a_750_n1638# a_n1954_n1768# 0.255f
C39 a_750_1206# a_n1954_n1768# 0.255f
C40 a_516_n1638# a_n1954_n1768# 0.255f
C41 a_516_1206# a_n1954_n1768# 0.255f
C42 a_282_n1638# a_n1954_n1768# 0.255f
C43 a_282_1206# a_n1954_n1768# 0.255f
C44 a_48_n1638# a_n1954_n1768# 0.255f
C45 a_48_1206# a_n1954_n1768# 0.255f
C46 a_n186_n1638# a_n1954_n1768# 0.255f
C47 a_n186_1206# a_n1954_n1768# 0.255f
C48 a_n420_n1638# a_n1954_n1768# 0.255f
C49 a_n420_1206# a_n1954_n1768# 0.255f
C50 a_n654_n1638# a_n1954_n1768# 0.255f
C51 a_n654_1206# a_n1954_n1768# 0.255f
C52 a_n888_n1638# a_n1954_n1768# 0.255f
C53 a_n888_1206# a_n1954_n1768# 0.255f
C54 a_n1122_n1638# a_n1954_n1768# 0.255f
C55 a_n1122_1206# a_n1954_n1768# 0.255f
C56 a_n1356_n1638# a_n1954_n1768# 0.255f
C57 a_n1356_1206# a_n1954_n1768# 0.255f
C58 a_n1590_n1638# a_n1954_n1768# 0.255f
C59 a_n1590_1206# a_n1954_n1768# 0.255f
C60 a_n1824_n1638# a_n1954_n1768# 0.465f
C61 a_n1824_1206# a_n1954_n1768# 0.465f
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_727CUP a_n100_n565# a_100_n477# a_n292_n699#
+ a_n158_n477#
X0 a_100_n477# a_n100_n565# a_n158_n477# a_n292_n699# sky130_fd_pr__nfet_g5v0d10v5 ad=1.38 pd=10.1 as=1.38 ps=10.1 w=4.77 l=1
C0 a_n158_n477# a_100_n477# 0.261f
C1 a_n100_n565# a_100_n477# 0.107f
C2 a_n100_n565# a_n158_n477# 0.107f
C3 a_100_n477# a_n292_n699# 0.53f
C4 a_n158_n477# a_n292_n699# 0.53f
C5 a_n100_n565# a_n292_n699# 0.714f
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_VU5C5A a_n287_n487# a_n421_n709# a_n229_n575#
+ a_229_n487# a_n29_n487# a_29_n575#
X0 a_229_n487# a_29_n575# a_n29_n487# a_n421_n709# sky130_fd_pr__nfet_g5v0d10v5 ad=1.41 pd=10.3 as=0.706 ps=5.16 w=4.87 l=1
X1 a_n29_n487# a_n229_n575# a_n287_n487# a_n421_n709# sky130_fd_pr__nfet_g5v0d10v5 ad=0.706 pd=5.16 as=1.41 ps=10.3 w=4.87 l=1
C0 a_n287_n487# a_n29_n487# 0.267f
C1 a_29_n575# a_n29_n487# 0.11f
C2 a_229_n487# a_n29_n487# 0.267f
C3 a_229_n487# a_29_n575# 0.11f
C4 a_n229_n575# a_n29_n487# 0.11f
C5 a_n229_n575# a_n287_n487# 0.11f
C6 a_n229_n575# a_29_n575# 0.104f
C7 a_229_n487# a_n421_n709# 0.54f
C8 a_n29_n487# a_n421_n709# 0.163f
C9 a_n287_n487# a_n421_n709# 0.54f
C10 a_29_n575# a_n421_n709# 0.651f
C11 a_n229_n575# a_n421_n709# 0.651f
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_J97EKB a_487_n438# a_n803_n438# a_29_n526# a_n745_n526#
+ a_n287_n438# a_n1061_n438# a_803_n526# a_745_n438# a_n229_n526# a_287_n526# a_n1003_n526#
+ a_229_n438# a_n545_n438# a_1003_n438# a_n487_n526# a_n1195_n660# a_545_n526# a_n29_n438#
X0 a_1003_n438# a_803_n526# a_745_n438# a_n1195_n660# sky130_fd_pr__nfet_g5v0d10v5 ad=1.27 pd=9.34 as=0.635 ps=4.67 w=4.38 l=1
X1 a_745_n438# a_545_n526# a_487_n438# a_n1195_n660# sky130_fd_pr__nfet_g5v0d10v5 ad=0.635 pd=4.67 as=0.635 ps=4.67 w=4.38 l=1
X2 a_487_n438# a_287_n526# a_229_n438# a_n1195_n660# sky130_fd_pr__nfet_g5v0d10v5 ad=0.635 pd=4.67 as=0.635 ps=4.67 w=4.38 l=1
X3 a_229_n438# a_29_n526# a_n29_n438# a_n1195_n660# sky130_fd_pr__nfet_g5v0d10v5 ad=0.635 pd=4.67 as=0.635 ps=4.67 w=4.38 l=1
X4 a_n29_n438# a_n229_n526# a_n287_n438# a_n1195_n660# sky130_fd_pr__nfet_g5v0d10v5 ad=0.635 pd=4.67 as=0.635 ps=4.67 w=4.38 l=1
X5 a_n545_n438# a_n745_n526# a_n803_n438# a_n1195_n660# sky130_fd_pr__nfet_g5v0d10v5 ad=0.635 pd=4.67 as=0.635 ps=4.67 w=4.38 l=1
X6 a_n287_n438# a_n487_n526# a_n545_n438# a_n1195_n660# sky130_fd_pr__nfet_g5v0d10v5 ad=0.635 pd=4.67 as=0.635 ps=4.67 w=4.38 l=1
X7 a_n803_n438# a_n1003_n526# a_n1061_n438# a_n1195_n660# sky130_fd_pr__nfet_g5v0d10v5 ad=0.635 pd=4.67 as=1.27 ps=9.34 w=4.38 l=1
C0 a_n545_n438# a_n487_n526# 0.099f
C1 a_n545_n438# a_n745_n526# 0.099f
C2 a_n803_n438# a_n745_n526# 0.099f
C3 a_229_n438# a_487_n438# 0.24f
C4 a_487_n438# a_745_n438# 0.24f
C5 a_745_n438# a_1003_n438# 0.24f
C6 a_n29_n438# a_229_n438# 0.24f
C7 a_n803_n438# a_n1061_n438# 0.24f
C8 a_n487_n526# a_n229_n526# 0.104f
C9 a_n745_n526# a_n487_n526# 0.104f
C10 a_29_n526# a_n229_n526# 0.104f
C11 a_487_n438# a_545_n526# 0.099f
C12 a_545_n526# a_745_n438# 0.099f
C13 a_29_n526# a_287_n526# 0.104f
C14 a_n29_n438# a_n287_n438# 0.24f
C15 a_n803_n438# a_n1003_n526# 0.099f
C16 a_n29_n438# a_n229_n526# 0.099f
C17 a_287_n526# a_487_n438# 0.099f
C18 a_287_n526# a_229_n438# 0.099f
C19 a_29_n526# a_229_n438# 0.099f
C20 a_29_n526# a_n29_n438# 0.099f
C21 a_803_n526# a_1003_n438# 0.099f
C22 a_n1003_n526# a_n745_n526# 0.104f
C23 a_803_n526# a_745_n438# 0.099f
C24 a_n545_n438# a_n287_n438# 0.24f
C25 a_n803_n438# a_n545_n438# 0.24f
C26 a_287_n526# a_545_n526# 0.104f
C27 a_n1061_n438# a_n1003_n526# 0.099f
C28 a_803_n526# a_545_n526# 0.104f
C29 a_n287_n438# a_n229_n526# 0.099f
C30 a_n287_n438# a_n487_n526# 0.099f
C31 a_1003_n438# a_n1195_n660# 0.489f
C32 a_745_n438# a_n1195_n660# 0.149f
C33 a_487_n438# a_n1195_n660# 0.149f
C34 a_229_n438# a_n1195_n660# 0.149f
C35 a_n29_n438# a_n1195_n660# 0.149f
C36 a_n287_n438# a_n1195_n660# 0.149f
C37 a_n545_n438# a_n1195_n660# 0.149f
C38 a_n803_n438# a_n1195_n660# 0.149f
C39 a_n1061_n438# a_n1195_n660# 0.489f
C40 a_803_n526# a_n1195_n660# 0.65f
C41 a_545_n526# a_n1195_n660# 0.587f
C42 a_287_n526# a_n1195_n660# 0.587f
C43 a_29_n526# a_n1195_n660# 0.587f
C44 a_n229_n526# a_n1195_n660# 0.587f
C45 a_n487_n526# a_n1195_n660# 0.587f
C46 a_n745_n526# a_n1195_n660# 0.587f
C47 a_n1003_n526# a_n1195_n660# 0.65f
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_S7E57E a_n229_n553# a_287_n553# a_229_n465# a_n545_n465#
+ a_n487_n553# a_487_n465# a_n29_n465# a_n679_n687# a_29_n553# a_n287_n465#
X0 a_487_n465# a_287_n553# a_229_n465# a_n679_n687# sky130_fd_pr__nfet_g5v0d10v5 ad=1.35 pd=9.88 as=0.674 ps=4.94 w=4.65 l=1
X1 a_229_n465# a_29_n553# a_n29_n465# a_n679_n687# sky130_fd_pr__nfet_g5v0d10v5 ad=0.674 pd=4.94 as=0.674 ps=4.94 w=4.65 l=1
X2 a_n29_n465# a_n229_n553# a_n287_n465# a_n679_n687# sky130_fd_pr__nfet_g5v0d10v5 ad=0.674 pd=4.94 as=0.674 ps=4.94 w=4.65 l=1
X3 a_n287_n465# a_n487_n553# a_n545_n465# a_n679_n687# sky130_fd_pr__nfet_g5v0d10v5 ad=0.674 pd=4.94 as=1.35 ps=9.88 w=4.65 l=1
C0 a_287_n553# a_229_n465# 0.105f
C1 a_29_n553# a_229_n465# 0.105f
C2 a_29_n553# a_287_n553# 0.104f
C3 a_n545_n465# a_n287_n465# 0.255f
C4 a_n229_n553# a_n287_n465# 0.105f
C5 a_n229_n553# a_29_n553# 0.104f
C6 a_n487_n553# a_n287_n465# 0.105f
C7 a_n487_n553# a_n545_n465# 0.105f
C8 a_n29_n465# a_229_n465# 0.255f
C9 a_n229_n553# a_n487_n553# 0.104f
C10 a_n29_n465# a_n287_n465# 0.255f
C11 a_29_n553# a_n29_n465# 0.105f
C12 a_n229_n553# a_n29_n465# 0.105f
C13 a_487_n465# a_229_n465# 0.255f
C14 a_287_n553# a_487_n465# 0.105f
C15 a_487_n465# a_n679_n687# 0.517f
C16 a_229_n465# a_n679_n687# 0.157f
C17 a_n29_n465# a_n679_n687# 0.157f
C18 a_n287_n465# a_n679_n687# 0.157f
C19 a_n545_n465# a_n679_n687# 0.517f
C20 a_287_n553# a_n679_n687# 0.651f
C21 a_29_n553# a_n679_n687# 0.588f
C22 a_n229_n553# a_n679_n687# 0.588f
C23 a_n487_n553# a_n679_n687# 0.651f
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_YPGNM4 a_545_n528# a_n545_n440# a_1577_n528#
+ a_1003_n440# a_n29_n440# a_29_n528# a_n1777_n528# a_487_n440# a_n745_n528# a_n1835_n440#
+ a_803_n528# a_n803_n440# a_1519_n440# a_1261_n440# a_n229_n528# a_n1319_n440# a_287_n528#
+ a_n1003_n528# a_n287_n440# a_n1061_n440# a_n1969_n662# a_745_n440# a_1319_n528#
+ a_1061_n528# a_1777_n440# a_n1519_n528# a_229_n440# a_n487_n528# a_n1261_n528# a_n1577_n440#
X0 a_1777_n440# a_1577_n528# a_1519_n440# a_n1969_n662# sky130_fd_pr__nfet_g5v0d10v5 ad=1.28 pd=9.38 as=0.638 ps=4.69 w=4.4 l=1
X1 a_1261_n440# a_1061_n528# a_1003_n440# a_n1969_n662# sky130_fd_pr__nfet_g5v0d10v5 ad=0.638 pd=4.69 as=0.638 ps=4.69 w=4.4 l=1
X2 a_229_n440# a_29_n528# a_n29_n440# a_n1969_n662# sky130_fd_pr__nfet_g5v0d10v5 ad=0.638 pd=4.69 as=0.638 ps=4.69 w=4.4 l=1
X3 a_n29_n440# a_n229_n528# a_n287_n440# a_n1969_n662# sky130_fd_pr__nfet_g5v0d10v5 ad=0.638 pd=4.69 as=0.638 ps=4.69 w=4.4 l=1
X4 a_n1319_n440# a_n1519_n528# a_n1577_n440# a_n1969_n662# sky130_fd_pr__nfet_g5v0d10v5 ad=0.638 pd=4.69 as=0.638 ps=4.69 w=4.4 l=1
X5 a_n545_n440# a_n745_n528# a_n803_n440# a_n1969_n662# sky130_fd_pr__nfet_g5v0d10v5 ad=0.638 pd=4.69 as=0.638 ps=4.69 w=4.4 l=1
X6 a_n803_n440# a_n1003_n528# a_n1061_n440# a_n1969_n662# sky130_fd_pr__nfet_g5v0d10v5 ad=0.638 pd=4.69 as=0.638 ps=4.69 w=4.4 l=1
X7 a_n287_n440# a_n487_n528# a_n545_n440# a_n1969_n662# sky130_fd_pr__nfet_g5v0d10v5 ad=0.638 pd=4.69 as=0.638 ps=4.69 w=4.4 l=1
X8 a_n1577_n440# a_n1777_n528# a_n1835_n440# a_n1969_n662# sky130_fd_pr__nfet_g5v0d10v5 ad=0.638 pd=4.69 as=1.28 ps=9.38 w=4.4 l=1
X9 a_1519_n440# a_1319_n528# a_1261_n440# a_n1969_n662# sky130_fd_pr__nfet_g5v0d10v5 ad=0.638 pd=4.69 as=0.638 ps=4.69 w=4.4 l=1
X10 a_n1061_n440# a_n1261_n528# a_n1319_n440# a_n1969_n662# sky130_fd_pr__nfet_g5v0d10v5 ad=0.638 pd=4.69 as=0.638 ps=4.69 w=4.4 l=1
X11 a_1003_n440# a_803_n528# a_745_n440# a_n1969_n662# sky130_fd_pr__nfet_g5v0d10v5 ad=0.638 pd=4.69 as=0.638 ps=4.69 w=4.4 l=1
X12 a_487_n440# a_287_n528# a_229_n440# a_n1969_n662# sky130_fd_pr__nfet_g5v0d10v5 ad=0.638 pd=4.69 as=0.638 ps=4.69 w=4.4 l=1
X13 a_745_n440# a_545_n528# a_487_n440# a_n1969_n662# sky130_fd_pr__nfet_g5v0d10v5 ad=0.638 pd=4.69 as=0.638 ps=4.69 w=4.4 l=1
C0 a_n1061_n440# a_n1003_n528# 0.0995f
C1 a_545_n528# a_803_n528# 0.104f
C2 a_n803_n440# a_n1003_n528# 0.0995f
C3 a_n1777_n528# a_n1519_n528# 0.104f
C4 a_n1519_n528# a_n1261_n528# 0.104f
C5 a_229_n440# a_487_n440# 0.241f
C6 a_n29_n440# a_229_n440# 0.241f
C7 a_545_n528# a_487_n440# 0.0995f
C8 a_n287_n440# a_n29_n440# 0.241f
C9 a_1003_n440# a_1261_n440# 0.241f
C10 a_287_n528# a_487_n440# 0.0995f
C11 a_287_n528# a_229_n440# 0.0995f
C12 a_745_n440# a_1003_n440# 0.241f
C13 a_n545_n440# a_n287_n440# 0.241f
C14 a_n1319_n440# a_n1061_n440# 0.241f
C15 a_n803_n440# a_n1061_n440# 0.241f
C16 a_n803_n440# a_n545_n440# 0.241f
C17 a_n1577_n440# a_n1319_n440# 0.241f
C18 a_n1777_n528# a_n1835_n440# 0.0995f
C19 a_287_n528# a_545_n528# 0.104f
C20 a_n229_n528# a_n29_n440# 0.0995f
C21 a_n287_n440# a_n229_n528# 0.0995f
C22 a_1261_n440# a_1319_n528# 0.0995f
C23 a_n287_n440# a_n487_n528# 0.0995f
C24 a_1519_n440# a_1777_n440# 0.241f
C25 a_n545_n440# a_n487_n528# 0.0995f
C26 a_n1003_n528# a_n745_n528# 0.104f
C27 a_n1003_n528# a_n1261_n528# 0.104f
C28 a_1261_n440# a_1061_n528# 0.0995f
C29 a_n487_n528# a_n229_n528# 0.104f
C30 a_1003_n440# a_1061_n528# 0.0995f
C31 a_1003_n440# a_803_n528# 0.0995f
C32 a_1319_n528# a_1577_n528# 0.104f
C33 a_745_n440# a_803_n528# 0.0995f
C34 a_29_n528# a_229_n440# 0.0995f
C35 a_29_n528# a_n29_n440# 0.0995f
C36 a_n545_n440# a_n745_n528# 0.0995f
C37 a_n1061_n440# a_n1261_n528# 0.0995f
C38 a_n803_n440# a_n745_n528# 0.0995f
C39 a_745_n440# a_487_n440# 0.241f
C40 a_n1319_n440# a_n1261_n528# 0.0995f
C41 a_1319_n528# a_1061_n528# 0.104f
C42 a_n1577_n440# a_n1777_n528# 0.0995f
C43 a_n1319_n440# a_n1519_n528# 0.0995f
C44 a_n1577_n440# a_n1519_n528# 0.0995f
C45 a_287_n528# a_29_n528# 0.104f
C46 a_545_n528# a_745_n440# 0.0995f
C47 a_1261_n440# a_1519_n440# 0.241f
C48 a_n487_n528# a_n745_n528# 0.104f
C49 a_29_n528# a_n229_n528# 0.104f
C50 a_803_n528# a_1061_n528# 0.104f
C51 a_n1577_n440# a_n1835_n440# 0.241f
C52 a_1777_n440# a_1577_n528# 0.0995f
C53 a_1519_n440# a_1577_n528# 0.0995f
C54 a_1519_n440# a_1319_n528# 0.0995f
C55 a_1777_n440# a_n1969_n662# 0.491f
C56 a_1519_n440# a_n1969_n662# 0.15f
C57 a_1261_n440# a_n1969_n662# 0.15f
C58 a_1003_n440# a_n1969_n662# 0.15f
C59 a_745_n440# a_n1969_n662# 0.15f
C60 a_487_n440# a_n1969_n662# 0.15f
C61 a_229_n440# a_n1969_n662# 0.15f
C62 a_n29_n440# a_n1969_n662# 0.15f
C63 a_n287_n440# a_n1969_n662# 0.15f
C64 a_n545_n440# a_n1969_n662# 0.15f
C65 a_n803_n440# a_n1969_n662# 0.15f
C66 a_n1061_n440# a_n1969_n662# 0.15f
C67 a_n1319_n440# a_n1969_n662# 0.15f
C68 a_n1577_n440# a_n1969_n662# 0.15f
C69 a_n1835_n440# a_n1969_n662# 0.491f
C70 a_1577_n528# a_n1969_n662# 0.65f
C71 a_1319_n528# a_n1969_n662# 0.587f
C72 a_1061_n528# a_n1969_n662# 0.587f
C73 a_803_n528# a_n1969_n662# 0.587f
C74 a_545_n528# a_n1969_n662# 0.587f
C75 a_287_n528# a_n1969_n662# 0.587f
C76 a_29_n528# a_n1969_n662# 0.587f
C77 a_n229_n528# a_n1969_n662# 0.587f
C78 a_n487_n528# a_n1969_n662# 0.587f
C79 a_n745_n528# a_n1969_n662# 0.587f
C80 a_n1003_n528# a_n1969_n662# 0.587f
C81 a_n1261_n528# a_n1969_n662# 0.587f
C82 a_n1519_n528# a_n1969_n662# 0.587f
C83 a_n1777_n528# a_n1969_n662# 0.65f
.ends

.subckt RB_array_20 VDD VSS R1 R2 D0 D1 D2 D3 D4
XXR1 VSS R2 m1_2651_1472# sky130_fd_pr__res_high_po_0p69_JKKHRG
XXR2 VSS R2 m1_2124_1470# sky130_fd_pr__res_high_po_0p69_JKKHRG
XXR3 R2 m1_3160_410# R2 VSS m1_3160_410# sky130_fd_pr__res_high_po_0p69_Z3RMRJ
XXR5 m1_5470_410# R2 R2 R2 m1_5470_410# R2 R2 m1_5470_410# R2 m1_5470_410# m1_5470_410#
+ m1_5470_410# m1_5470_410# R2 VSS R2 m1_5470_410# sky130_fd_pr__res_high_po_0p69_Z3RMR6
XXR4 R2 VSS m1_4060_410# R2 R2 m1_4060_410# m1_4060_410# m1_4060_410# R2 sky130_fd_pr__res_high_po_0p69_YMHKRJ
XXR6 m1_7940_410# R2 R2 R2 R2 m1_7940_410# m1_7940_410# m1_7940_410# R2 VSS R2 R2
+ m1_7940_410# R2 m1_7940_410# R2 R2 m1_7940_410# m1_7940_410# R2 R2 R2 m1_7940_410#
+ m1_7940_410# m1_7940_410# m1_7940_410# R2 R2 m1_7940_410# m1_7940_410# R2 m1_7940_410#
+ m1_7940_410# sky130_fd_pr__res_high_po_0p69_HBQF5Z
XXM6 D0 m1_2651_1472# VSS R1 sky130_fd_pr__nfet_g5v0d10v5_727CUP
XXM7 m1_3160_410# VSS D1 m1_3160_410# R1 D1 sky130_fd_pr__nfet_g5v0d10v5_VU5C5A
XXM9 m1_5470_410# R1 D3 D3 R1 m1_5470_410# D3 R1 D3 D3 D3 R1 m1_5470_410# m1_5470_410#
+ D3 VSS D3 m1_5470_410# sky130_fd_pr__nfet_g5v0d10v5_J97EKB
XXM8 D2 D2 R1 m1_4060_410# D2 m1_4060_410# m1_4060_410# VSS D2 R1 sky130_fd_pr__nfet_g5v0d10v5_S7E57E
XXM10 D4 R1 D4 R1 R1 D4 D4 R1 D4 m1_7940_410# D4 m1_7940_410# R1 m1_7940_410# D4 m1_7940_410#
+ D4 D4 m1_7940_410# R1 VSS m1_7940_410# D4 D4 m1_7940_410# D4 m1_7940_410# D4 D4
+ R1 sky130_fd_pr__nfet_g5v0d10v5_YPGNM4
XXM11 VDD m1_2124_1470# VSS R1 sky130_fd_pr__nfet_g5v0d10v5_727CUP
C0 m1_2651_1472# D0 0.449f
C1 m1_2651_1472# D3 0.0446f
C2 D4 m1_3160_410# 0.458f
C3 D1 m1_2124_1470# 0.0674f
C4 D0 R1 0.619f
C5 R1 D3 4.08f
C6 D0 VDD 0.332f
C7 m1_3160_410# m1_4060_410# 0.201f
C8 D2 m1_3160_410# 0.163f
C9 D3 VDD 0.0728f
C10 D3 m1_5470_410# 3.93f
C11 m1_2651_1472# R1 -0.107f
C12 D1 m1_3160_410# 1.09f
C13 D0 D4 0.0964f
C14 D3 D4 3.99f
C15 D0 m1_4060_410# 7.28e-21
C16 D0 D2 0.0732f
C17 m1_3160_410# m1_2124_1470# 1.43e-19
C18 R1 VDD 0.551f
C19 D3 m1_4060_410# 0.2f
C20 D2 D3 2.27f
C21 D3 m1_7940_410# 5.93e-19
C22 R1 m1_5470_410# 0.379f
C23 m1_2651_1472# D4 0.0516f
C24 D0 D1 0.731f
C25 m1_2651_1472# m1_4060_410# 2.22e-21
C26 D3 D1 0.145f
C27 m1_2651_1472# D2 0.0483f
C28 R1 D4 7.57f
C29 VDD D4 0.0966f
C30 D0 m1_2124_1470# 0.126f
C31 R1 m1_4060_410# 0.226f
C32 D2 R1 2.15f
C33 D3 m1_2124_1470# 0.0433f
C34 D2 VDD 0.0734f
C35 D4 m1_5470_410# 1.37f
C36 R1 m1_7940_410# 0.29f
C37 m1_2651_1472# D1 0.114f
C38 m1_4060_410# m1_5470_410# 0.176f
C39 D2 m1_5470_410# 5.82e-19
C40 R1 D1 1.16f
C41 m1_7940_410# m1_5470_410# 0.197f
C42 m1_2651_1472# m1_2124_1470# 0.104f
C43 VDD D1 0.0754f
C44 D0 m1_3160_410# 0.00189f
C45 D4 m1_4060_410# 0.742f
C46 D2 D4 0.308f
C47 D3 m1_3160_410# 0.12f
C48 R1 m1_2124_1470# 0.0621f
C49 D4 m1_7940_410# 8.65f
C50 D2 m1_4060_410# 2.08f
C51 VDD m1_2124_1470# 0.494f
C52 D4 D1 0.154f
C53 m1_2651_1472# m1_3160_410# 0.19f
C54 D1 m1_4060_410# 1.86e-19
C55 D2 D1 1.31f
C56 D4 m1_2124_1470# 0.0503f
C57 R1 m1_3160_410# 0.177f
C58 D0 D3 0.0725f
C59 VDD m1_3160_410# 4.48e-19
C60 D2 m1_2124_1470# 0.0469f
C61 R1 VSS 4.54f
C62 VDD VSS 0.914f
C63 m1_7940_410# VSS 7.18f
C64 D4 VSS 8.99f
C65 D2 VSS 2.7f
C66 D3 VSS 5.24f
C67 D1 VSS 1.48f
C68 D0 VSS 0.884f
C69 m1_4060_410# VSS 3.17f
C70 m1_5470_410# VSS 4.68f
C71 m1_3160_410# VSS 2.43f
C72 R2 VSS 15.3f
C73 m1_2124_1470# VSS 1.55f
C74 m1_2651_1472# VSS 1.58f
.ends

