magic
tech sky130A
magscale 1 2
timestamp 1718246682
<< pwell >>
rect -1231 -696 1231 696
<< mvnmos >>
rect -1003 -438 -803 438
rect -745 -438 -545 438
rect -487 -438 -287 438
rect -229 -438 -29 438
rect 29 -438 229 438
rect 287 -438 487 438
rect 545 -438 745 438
rect 803 -438 1003 438
<< mvndiff >>
rect -1061 426 -1003 438
rect -1061 -426 -1049 426
rect -1015 -426 -1003 426
rect -1061 -438 -1003 -426
rect -803 426 -745 438
rect -803 -426 -791 426
rect -757 -426 -745 426
rect -803 -438 -745 -426
rect -545 426 -487 438
rect -545 -426 -533 426
rect -499 -426 -487 426
rect -545 -438 -487 -426
rect -287 426 -229 438
rect -287 -426 -275 426
rect -241 -426 -229 426
rect -287 -438 -229 -426
rect -29 426 29 438
rect -29 -426 -17 426
rect 17 -426 29 426
rect -29 -438 29 -426
rect 229 426 287 438
rect 229 -426 241 426
rect 275 -426 287 426
rect 229 -438 287 -426
rect 487 426 545 438
rect 487 -426 499 426
rect 533 -426 545 426
rect 487 -438 545 -426
rect 745 426 803 438
rect 745 -426 757 426
rect 791 -426 803 426
rect 745 -438 803 -426
rect 1003 426 1061 438
rect 1003 -426 1015 426
rect 1049 -426 1061 426
rect 1003 -438 1061 -426
<< mvndiffc >>
rect -1049 -426 -1015 426
rect -791 -426 -757 426
rect -533 -426 -499 426
rect -275 -426 -241 426
rect -17 -426 17 426
rect 241 -426 275 426
rect 499 -426 533 426
rect 757 -426 791 426
rect 1015 -426 1049 426
<< mvpsubdiff >>
rect -1195 648 1195 660
rect -1195 614 -1087 648
rect 1087 614 1195 648
rect -1195 602 1195 614
rect -1195 552 -1137 602
rect -1195 -552 -1183 552
rect -1149 -552 -1137 552
rect 1137 552 1195 602
rect -1195 -602 -1137 -552
rect 1137 -552 1149 552
rect 1183 -552 1195 552
rect 1137 -602 1195 -552
rect -1195 -614 1195 -602
rect -1195 -648 -1087 -614
rect 1087 -648 1195 -614
rect -1195 -660 1195 -648
<< mvpsubdiffcont >>
rect -1087 614 1087 648
rect -1183 -552 -1149 552
rect 1149 -552 1183 552
rect -1087 -648 1087 -614
<< poly >>
rect -1003 510 -803 526
rect -1003 476 -987 510
rect -819 476 -803 510
rect -1003 438 -803 476
rect -745 510 -545 526
rect -745 476 -729 510
rect -561 476 -545 510
rect -745 438 -545 476
rect -487 510 -287 526
rect -487 476 -471 510
rect -303 476 -287 510
rect -487 438 -287 476
rect -229 510 -29 526
rect -229 476 -213 510
rect -45 476 -29 510
rect -229 438 -29 476
rect 29 510 229 526
rect 29 476 45 510
rect 213 476 229 510
rect 29 438 229 476
rect 287 510 487 526
rect 287 476 303 510
rect 471 476 487 510
rect 287 438 487 476
rect 545 510 745 526
rect 545 476 561 510
rect 729 476 745 510
rect 545 438 745 476
rect 803 510 1003 526
rect 803 476 819 510
rect 987 476 1003 510
rect 803 438 1003 476
rect -1003 -476 -803 -438
rect -1003 -510 -987 -476
rect -819 -510 -803 -476
rect -1003 -526 -803 -510
rect -745 -476 -545 -438
rect -745 -510 -729 -476
rect -561 -510 -545 -476
rect -745 -526 -545 -510
rect -487 -476 -287 -438
rect -487 -510 -471 -476
rect -303 -510 -287 -476
rect -487 -526 -287 -510
rect -229 -476 -29 -438
rect -229 -510 -213 -476
rect -45 -510 -29 -476
rect -229 -526 -29 -510
rect 29 -476 229 -438
rect 29 -510 45 -476
rect 213 -510 229 -476
rect 29 -526 229 -510
rect 287 -476 487 -438
rect 287 -510 303 -476
rect 471 -510 487 -476
rect 287 -526 487 -510
rect 545 -476 745 -438
rect 545 -510 561 -476
rect 729 -510 745 -476
rect 545 -526 745 -510
rect 803 -476 1003 -438
rect 803 -510 819 -476
rect 987 -510 1003 -476
rect 803 -526 1003 -510
<< polycont >>
rect -987 476 -819 510
rect -729 476 -561 510
rect -471 476 -303 510
rect -213 476 -45 510
rect 45 476 213 510
rect 303 476 471 510
rect 561 476 729 510
rect 819 476 987 510
rect -987 -510 -819 -476
rect -729 -510 -561 -476
rect -471 -510 -303 -476
rect -213 -510 -45 -476
rect 45 -510 213 -476
rect 303 -510 471 -476
rect 561 -510 729 -476
rect 819 -510 987 -476
<< locali >>
rect -1183 614 -1087 648
rect 1087 614 1183 648
rect -1183 552 -1149 614
rect 1149 552 1183 614
rect -1003 476 -987 510
rect -819 476 -803 510
rect -745 476 -729 510
rect -561 476 -545 510
rect -487 476 -471 510
rect -303 476 -287 510
rect -229 476 -213 510
rect -45 476 -29 510
rect 29 476 45 510
rect 213 476 229 510
rect 287 476 303 510
rect 471 476 487 510
rect 545 476 561 510
rect 729 476 745 510
rect 803 476 819 510
rect 987 476 1003 510
rect -1049 426 -1015 442
rect -1049 -442 -1015 -426
rect -791 426 -757 442
rect -791 -442 -757 -426
rect -533 426 -499 442
rect -533 -442 -499 -426
rect -275 426 -241 442
rect -275 -442 -241 -426
rect -17 426 17 442
rect -17 -442 17 -426
rect 241 426 275 442
rect 241 -442 275 -426
rect 499 426 533 442
rect 499 -442 533 -426
rect 757 426 791 442
rect 757 -442 791 -426
rect 1015 426 1049 442
rect 1015 -442 1049 -426
rect -1003 -510 -987 -476
rect -819 -510 -803 -476
rect -745 -510 -729 -476
rect -561 -510 -545 -476
rect -487 -510 -471 -476
rect -303 -510 -287 -476
rect -229 -510 -213 -476
rect -45 -510 -29 -476
rect 29 -510 45 -476
rect 213 -510 229 -476
rect 287 -510 303 -476
rect 471 -510 487 -476
rect 545 -510 561 -476
rect 729 -510 745 -476
rect 803 -510 819 -476
rect 987 -510 1003 -476
rect -1183 -614 -1149 -552
rect 1149 -614 1183 -552
rect -1183 -648 -1087 -614
rect 1087 -648 1183 -614
<< viali >>
rect -987 476 -819 510
rect -729 476 -561 510
rect -471 476 -303 510
rect -213 476 -45 510
rect 45 476 213 510
rect 303 476 471 510
rect 561 476 729 510
rect 819 476 987 510
rect -1049 -426 -1015 426
rect -791 -426 -757 426
rect -533 -426 -499 426
rect -275 -426 -241 426
rect -17 -426 17 426
rect 241 -426 275 426
rect 499 -426 533 426
rect 757 -426 791 426
rect 1015 -426 1049 426
rect -987 -510 -819 -476
rect -729 -510 -561 -476
rect -471 -510 -303 -476
rect -213 -510 -45 -476
rect 45 -510 213 -476
rect 303 -510 471 -476
rect 561 -510 729 -476
rect 819 -510 987 -476
<< metal1 >>
rect -999 510 -807 516
rect -999 476 -987 510
rect -819 476 -807 510
rect -999 470 -807 476
rect -741 510 -549 516
rect -741 476 -729 510
rect -561 476 -549 510
rect -741 470 -549 476
rect -483 510 -291 516
rect -483 476 -471 510
rect -303 476 -291 510
rect -483 470 -291 476
rect -225 510 -33 516
rect -225 476 -213 510
rect -45 476 -33 510
rect -225 470 -33 476
rect 33 510 225 516
rect 33 476 45 510
rect 213 476 225 510
rect 33 470 225 476
rect 291 510 483 516
rect 291 476 303 510
rect 471 476 483 510
rect 291 470 483 476
rect 549 510 741 516
rect 549 476 561 510
rect 729 476 741 510
rect 549 470 741 476
rect 807 510 999 516
rect 807 476 819 510
rect 987 476 999 510
rect 807 470 999 476
rect -1055 426 -1009 438
rect -1055 -426 -1049 426
rect -1015 -426 -1009 426
rect -1055 -438 -1009 -426
rect -797 426 -751 438
rect -797 -426 -791 426
rect -757 -426 -751 426
rect -797 -438 -751 -426
rect -539 426 -493 438
rect -539 -426 -533 426
rect -499 -426 -493 426
rect -539 -438 -493 -426
rect -281 426 -235 438
rect -281 -426 -275 426
rect -241 -426 -235 426
rect -281 -438 -235 -426
rect -23 426 23 438
rect -23 -426 -17 426
rect 17 -426 23 426
rect -23 -438 23 -426
rect 235 426 281 438
rect 235 -426 241 426
rect 275 -426 281 426
rect 235 -438 281 -426
rect 493 426 539 438
rect 493 -426 499 426
rect 533 -426 539 426
rect 493 -438 539 -426
rect 751 426 797 438
rect 751 -426 757 426
rect 791 -426 797 426
rect 751 -438 797 -426
rect 1009 426 1055 438
rect 1009 -426 1015 426
rect 1049 -426 1055 426
rect 1009 -438 1055 -426
rect -999 -476 -807 -470
rect -999 -510 -987 -476
rect -819 -510 -807 -476
rect -999 -516 -807 -510
rect -741 -476 -549 -470
rect -741 -510 -729 -476
rect -561 -510 -549 -476
rect -741 -516 -549 -510
rect -483 -476 -291 -470
rect -483 -510 -471 -476
rect -303 -510 -291 -476
rect -483 -516 -291 -510
rect -225 -476 -33 -470
rect -225 -510 -213 -476
rect -45 -510 -33 -476
rect -225 -516 -33 -510
rect 33 -476 225 -470
rect 33 -510 45 -476
rect 213 -510 225 -476
rect 33 -516 225 -510
rect 291 -476 483 -470
rect 291 -510 303 -476
rect 471 -510 483 -476
rect 291 -516 483 -510
rect 549 -476 741 -470
rect 549 -510 561 -476
rect 729 -510 741 -476
rect 549 -516 741 -510
rect 807 -476 999 -470
rect 807 -510 819 -476
rect 987 -510 999 -476
rect 807 -516 999 -510
<< properties >>
string FIXED_BBOX -1166 -631 1166 631
string gencell sky130_fd_pr__nfet_g5v0d10v5
string library sky130
string parameters w 4.38 l 1.0 m 1 nf 8 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
