magic
tech sky130A
magscale 1 2
timestamp 1718246682
<< nwell >>
rect -745 -2197 745 2197
<< mvpmos >>
rect -487 -1900 -287 1900
rect -229 -1900 -29 1900
rect 29 -1900 229 1900
rect 287 -1900 487 1900
<< mvpdiff >>
rect -545 1888 -487 1900
rect -545 -1888 -533 1888
rect -499 -1888 -487 1888
rect -545 -1900 -487 -1888
rect -287 1888 -229 1900
rect -287 -1888 -275 1888
rect -241 -1888 -229 1888
rect -287 -1900 -229 -1888
rect -29 1888 29 1900
rect -29 -1888 -17 1888
rect 17 -1888 29 1888
rect -29 -1900 29 -1888
rect 229 1888 287 1900
rect 229 -1888 241 1888
rect 275 -1888 287 1888
rect 229 -1900 287 -1888
rect 487 1888 545 1900
rect 487 -1888 499 1888
rect 533 -1888 545 1888
rect 487 -1900 545 -1888
<< mvpdiffc >>
rect -533 -1888 -499 1888
rect -275 -1888 -241 1888
rect -17 -1888 17 1888
rect 241 -1888 275 1888
rect 499 -1888 533 1888
<< mvnsubdiff >>
rect -679 2119 679 2131
rect -679 2085 -571 2119
rect 571 2085 679 2119
rect -679 2073 679 2085
rect -679 2023 -621 2073
rect -679 -2023 -667 2023
rect -633 -2023 -621 2023
rect 621 2023 679 2073
rect -679 -2073 -621 -2023
rect 621 -2023 633 2023
rect 667 -2023 679 2023
rect 621 -2073 679 -2023
rect -679 -2085 679 -2073
rect -679 -2119 -571 -2085
rect 571 -2119 679 -2085
rect -679 -2131 679 -2119
<< mvnsubdiffcont >>
rect -571 2085 571 2119
rect -667 -2023 -633 2023
rect 633 -2023 667 2023
rect -571 -2119 571 -2085
<< poly >>
rect -487 1981 -287 1997
rect -487 1947 -471 1981
rect -303 1947 -287 1981
rect -487 1900 -287 1947
rect -229 1981 -29 1997
rect -229 1947 -213 1981
rect -45 1947 -29 1981
rect -229 1900 -29 1947
rect 29 1981 229 1997
rect 29 1947 45 1981
rect 213 1947 229 1981
rect 29 1900 229 1947
rect 287 1981 487 1997
rect 287 1947 303 1981
rect 471 1947 487 1981
rect 287 1900 487 1947
rect -487 -1947 -287 -1900
rect -487 -1981 -471 -1947
rect -303 -1981 -287 -1947
rect -487 -1997 -287 -1981
rect -229 -1947 -29 -1900
rect -229 -1981 -213 -1947
rect -45 -1981 -29 -1947
rect -229 -1997 -29 -1981
rect 29 -1947 229 -1900
rect 29 -1981 45 -1947
rect 213 -1981 229 -1947
rect 29 -1997 229 -1981
rect 287 -1947 487 -1900
rect 287 -1981 303 -1947
rect 471 -1981 487 -1947
rect 287 -1997 487 -1981
<< polycont >>
rect -471 1947 -303 1981
rect -213 1947 -45 1981
rect 45 1947 213 1981
rect 303 1947 471 1981
rect -471 -1981 -303 -1947
rect -213 -1981 -45 -1947
rect 45 -1981 213 -1947
rect 303 -1981 471 -1947
<< locali >>
rect -667 2085 -571 2119
rect 571 2085 667 2119
rect -667 2023 -633 2085
rect 633 2023 667 2085
rect -487 1947 -471 1981
rect -303 1947 -287 1981
rect -229 1947 -213 1981
rect -45 1947 -29 1981
rect 29 1947 45 1981
rect 213 1947 229 1981
rect 287 1947 303 1981
rect 471 1947 487 1981
rect -533 1888 -499 1904
rect -533 -1904 -499 -1888
rect -275 1888 -241 1904
rect -275 -1904 -241 -1888
rect -17 1888 17 1904
rect -17 -1904 17 -1888
rect 241 1888 275 1904
rect 241 -1904 275 -1888
rect 499 1888 533 1904
rect 499 -1904 533 -1888
rect -487 -1981 -471 -1947
rect -303 -1981 -287 -1947
rect -229 -1981 -213 -1947
rect -45 -1981 -29 -1947
rect 29 -1981 45 -1947
rect 213 -1981 229 -1947
rect 287 -1981 303 -1947
rect 471 -1981 487 -1947
rect -667 -2085 -633 -2023
rect 633 -2085 667 -2023
rect -667 -2119 -571 -2085
rect 571 -2119 667 -2085
<< viali >>
rect -471 1947 -303 1981
rect -213 1947 -45 1981
rect 45 1947 213 1981
rect 303 1947 471 1981
rect -533 -1888 -499 1888
rect -275 -1888 -241 1888
rect -17 -1888 17 1888
rect 241 -1888 275 1888
rect 499 -1888 533 1888
rect -471 -1981 -303 -1947
rect -213 -1981 -45 -1947
rect 45 -1981 213 -1947
rect 303 -1981 471 -1947
<< metal1 >>
rect -483 1981 -291 1987
rect -483 1947 -471 1981
rect -303 1947 -291 1981
rect -483 1941 -291 1947
rect -225 1981 -33 1987
rect -225 1947 -213 1981
rect -45 1947 -33 1981
rect -225 1941 -33 1947
rect 33 1981 225 1987
rect 33 1947 45 1981
rect 213 1947 225 1981
rect 33 1941 225 1947
rect 291 1981 483 1987
rect 291 1947 303 1981
rect 471 1947 483 1981
rect 291 1941 483 1947
rect -539 1888 -493 1900
rect -539 -1888 -533 1888
rect -499 -1888 -493 1888
rect -539 -1900 -493 -1888
rect -281 1888 -235 1900
rect -281 -1888 -275 1888
rect -241 -1888 -235 1888
rect -281 -1900 -235 -1888
rect -23 1888 23 1900
rect -23 -1888 -17 1888
rect 17 -1888 23 1888
rect -23 -1900 23 -1888
rect 235 1888 281 1900
rect 235 -1888 241 1888
rect 275 -1888 281 1888
rect 235 -1900 281 -1888
rect 493 1888 539 1900
rect 493 -1888 499 1888
rect 533 -1888 539 1888
rect 493 -1900 539 -1888
rect -483 -1947 -291 -1941
rect -483 -1981 -471 -1947
rect -303 -1981 -291 -1947
rect -483 -1987 -291 -1981
rect -225 -1947 -33 -1941
rect -225 -1981 -213 -1947
rect -45 -1981 -33 -1947
rect -225 -1987 -33 -1981
rect 33 -1947 225 -1941
rect 33 -1981 45 -1947
rect 213 -1981 225 -1947
rect 33 -1987 225 -1981
rect 291 -1947 483 -1941
rect 291 -1981 303 -1947
rect 471 -1981 483 -1947
rect 291 -1987 483 -1981
<< properties >>
string FIXED_BBOX -650 -2102 650 2102
string gencell sky130_fd_pr__pfet_g5v0d10v5
string library sky130
string parameters w 19.0 l 1.0 m 1 nf 4 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
