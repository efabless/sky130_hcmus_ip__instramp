* NGSPICE file created from sky130_hcmus_ip__instramp.ext - technology: sky130A

.subckt sky130_hcmus_ip__instramp AVOUT2 D5 V2 ibias G D0 D6 D2 D8 VSS AVOUT1 VOUT
+ V1 D1 D4 D3 ena D7 DVDD D9 VDD DVSS
X0 x6.V1.t40 x9.V2.t27 VSS.t160 sky130_fd_pr__res_high_po_0p69 l=12.22
X1 ia_opamp_0.V2.t37 a_1031_764.t4 VDD.t233 VDD.t232 sky130_fd_pr__pfet_g5v0d10v5 ad=2.755 pd=19.29 as=2.755 ps=19.29 w=19 l=1
X2 a_n2577_n5175# a_n2603_n5122# DVSS.t131 DVSS.t126 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X3 x6.V1.t18 D93v3.t2 a_16261_n9984.t27 VSS.t81 sky130_fd_pr__nfet_g5v0d10v5 ad=0.638 pd=4.69 as=0.638 ps=4.69 w=4.4 l=1
X4 VOUT.t33 a_16951_764.t4 VDD.t34 VDD.t33 sky130_fd_pr__pfet_g5v0d10v5 ad=2.755 pd=19.29 as=2.755 ps=19.29 w=19 l=1
X5 DVDD.t37 a_n2559_13399# a_n2603_12350# DVDD.t36 sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.12 as=0.2478 ps=2.27 w=0.84 l=0.15
X6 x6.V1.t79 x9.V2.t57 VSS.t199 sky130_fd_pr__res_high_po_0p69 l=12.22
X7 x3.R1.t79 D93v3.t3 a_16261_n4916.t27 VSS.t81 sky130_fd_pr__nfet_g5v0d10v5 ad=0.638 pd=4.69 as=0.638 ps=4.69 w=4.4 l=1
X8 DVSS.t214 a_n2559_3415# a_n2121_2781# DVSS.t213 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X9 x5.V2.t0 x4.V2.t0 VSS.t0 sky130_fd_pr__res_high_po_0p69 l=12.22
X10 DVSS.t87 a_n2559_n1577# a_n2121_n2211# DVSS.t86 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.3975 ps=3.53 w=1.5 l=0.5
X11 a_6164_n9984.t17 D43v3.t2 x5.V2.t47 VSS.t18 sky130_fd_pr__nfet_g5v0d10v5 ad=0.638 pd=4.69 as=0.638 ps=4.69 w=4.4 l=1
X12 AVOUT2.t29 a_6164_n9984.t25 VSS.t236 sky130_fd_pr__res_high_po_0p69 l=12.22
X13 x5.V2.t26 D33v3.t2 a_3720_n9984.t10 VSS.t124 sky130_fd_pr__nfet_g5v0d10v5 ad=0.6351 pd=4.67 as=1.2702 ps=9.34 w=4.38 l=1
X14 x6.V1.t80 x9.V2.t58 VSS.t0 sky130_fd_pr__res_high_po_0p69 l=12.22
X15 a_6164_n4916.t18 D43v3.t3 x4.V2.t5 VSS.t18 sky130_fd_pr__nfet_g5v0d10v5 ad=0.638 pd=4.69 as=0.638 ps=4.69 w=4.4 l=1
X16 AVOUT1.t32 a_6164_n4916.t27 VSS.t236 sky130_fd_pr__res_high_po_0p69 l=12.22
X17 x6.V1.t41 x9.V2.t28 VSS.t158 sky130_fd_pr__res_high_po_0p69 l=12.22
X18 x6.V1.t83 D73v3.t2 a_12405_n9984.t5 VSS.t75 sky130_fd_pr__nfet_g5v0d10v5 ad=0.67425 pd=4.94 as=1.3485 ps=9.88 w=4.65 l=1
X19 x4.V2.t60 D33v3.t3 a_3720_n4916.t9 VSS.t124 sky130_fd_pr__nfet_g5v0d10v5 ad=0.6351 pd=4.67 as=1.2702 ps=9.34 w=4.38 l=1
X20 x6.V1.t78 x9.V2.t56 VSS.t107 sky130_fd_pr__res_high_po_0p69 l=12.22
X21 x3.R1.t80 x8.V2.t57 VSS.t13 sky130_fd_pr__res_high_po_0p69 l=12.22
X22 x3.R1.t15 D73v3.t3 a_12405_n4916.t6 VSS.t75 sky130_fd_pr__nfet_g5v0d10v5 ad=0.67425 pd=4.94 as=1.3485 ps=9.88 w=4.65 l=1
X23 a_n2121_n4707# a_n2577_n5175# VDD.t110 VDD.t109 sky130_fd_pr__pfet_g5v0d10v5 ad=0.2142 pd=1.99 as=0.2142 ps=1.99 w=0.42 l=1
X24 DVDD.t25 a_n2559_15895# a_n2603_14846# DVDD.t24 sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.12 as=0.2478 ps=2.27 w=0.84 l=0.15
X25 x3.R1.t38 x8.V2.t37 VSS.t30 sky130_fd_pr__res_high_po_0p69 l=12.22
X26 ia_opamp_0.V2.t21 a_16261_n9984.t11 VSS.t148 sky130_fd_pr__res_high_po_0p69 l=12.22
X27 a_230_281.t0 ia_opamp_0.V2.t12 VSS.t139 sky130_fd_pr__res_high_po_0p69 l=3.2
X28 a_16951_764.t0 a_16157_764.t5 VDD.t3 VDD.t2 sky130_fd_pr__pfet_g5v0d10v5 ad=2.175 pd=15.29 as=4.35 ps=30.58 w=15 l=1
X29 a_6605_764.t3 a_6605_764.t2 VDD.t50 VDD.t49 sky130_fd_pr__pfet_g5v0d10v5 ad=2.175 pd=15.29 as=4.35 ps=30.58 w=15 l=1
X30 a_n2121_285# a_n2577_n183# VDD.t54 VDD.t53 sky130_fd_pr__pfet_g5v0d10v5 ad=0.2142 pd=1.99 as=0.2142 ps=1.99 w=0.42 l=1
X31 DVSS.t93 a_n2603_n7618# a_n2577_n7671# DVSS.t88 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X32 VOUT.t13 a_16261_n4916.t4 VSS.t148 sky130_fd_pr__res_high_po_0p69 l=12.22
X33 a_n2121_5277# a_n2559_5911# DVSS.t68 DVSS.t67 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X34 ia_opamp_0.V2.t20 a_13817_n9984.t4 VSS.t187 sky130_fd_pr__res_high_po_0p69 l=12.22
X35 a_n1825_n338# a_n2121_285# VDD.t57 VDD.t8 sky130_fd_pr__pfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.24375 ps=1.825 w=1.5 l=0.5
X36 a_n2577_14793# a_n2121_15261# VDD.t194 VDD.t193 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1365 pd=1.49 as=0.1113 ps=1.37 w=0.42 l=1
X37 DVSS.t85 a_n2559_n1577# a_n2603_n2626# DVSS.t84 sky130_fd_pr__nfet_01v8 ad=0.1176 pd=1.12 as=0.2478 ps=2.27 w=0.84 l=0.15
X38 x3.R1.t90 x8.V2.t67 VSS.t98 sky130_fd_pr__res_high_po_0p69 l=12.22
X39 VOUT.t37 a_13817_n4916.t15 VSS.t187 sky130_fd_pr__res_high_po_0p69 l=12.22
X40 DVSS.t111 D9.t0 sky130_fd_pr__diode_pw2nd_11v0 perim=3.16e+06 area=6.072e+11
X41 VDD.t156 DVSS.t307 VDD.t155 VDD.t154 sky130_fd_pr__pfet_g5v0d10v5 ad=0.265 pd=2.53 as=0 ps=0 w=1 l=1
X42 x3.R1.t86 x8.V2.t63 VSS.t177 sky130_fd_pr__res_high_po_0p69 l=12.22
X43 a_11509_n9984# D63v3.t2 x6.V1.t82 VSS.t220 sky130_fd_pr__nfet_g5v0d10v5 ad=1.4123 pd=10.32 as=0.70615 ps=5.16 w=4.87 l=1
X44 x6.V1.t57 x9.V2.t42 VSS.t13 sky130_fd_pr__res_high_po_0p69 l=12.22
X45 x5.V2.t6 x4.V2.t7 VSS.t29 sky130_fd_pr__res_high_po_0p69 l=12.22
X46 a_11509_n4916# D63v3.t3 x3.R1.t55 VSS.t220 sky130_fd_pr__nfet_g5v0d10v5 ad=1.4123 pd=10.32 as=0.70615 ps=5.16 w=4.87 l=1
X47 x5.V2.t38 x4.V2.t38 VSS.t94 sky130_fd_pr__res_high_po_0p69 l=12.22
X48 DVSS.t27 a_n2603_n10114# a_n2577_n10167# DVSS.t22 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X49 x6.V1.t8 x9.V2.t2 VSS.t30 sky130_fd_pr__res_high_po_0p69 l=12.22
X50 a_16150_281.t1 a_16951_764.t1 sky130_fd_pr__cap_mim_m3_1 l=6.9 w=6.9
X51 a_n2121_285# a_n2559_919# DVSS.t268 DVSS.t267 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X52 x5.V2.t5 D43v3.t4 a_6164_n9984.t16 VSS.t19 sky130_fd_pr__nfet_g5v0d10v5 ad=0.638 pd=4.69 as=0.638 ps=4.69 w=4.4 l=1
X53 x3.R1.t83 x8.V2.t60 VSS.t14 sky130_fd_pr__res_high_po_0p69 l=12.22
X54 AVOUT2.t11 a_1412_n9984# VSS.t41 sky130_fd_pr__res_high_po_0p69 l=12.22
X55 x4.V2.t6 D43v3.t5 a_6164_n4916.t17 VSS.t19 sky130_fd_pr__nfet_g5v0d10v5 ad=0.638 pd=4.69 as=0.638 ps=4.69 w=4.4 l=1
X56 AVOUT1.t5 a_1412_n4916# VSS.t41 sky130_fd_pr__res_high_po_0p69 l=12.22
X57 a_12973_764.t3 a_12973_764.t2 VDD.t134 VDD.t133 sky130_fd_pr__pfet_g5v0d10v5 ad=2.175 pd=15.29 as=4.35 ps=30.58 w=15 l=1
X58 x6.V1.t24 x9.V2.t12 VSS.t98 sky130_fd_pr__res_high_po_0p69 l=12.22
X59 x5.V2.t80 x4.V2.t81 VSS.t91 sky130_fd_pr__res_high_po_0p69 l=12.22
X60 ia_opamp_0.V2.t15 a_11509_n9984# VSS.t99 sky130_fd_pr__res_high_po_0p69 l=12.22
X61 AVOUT2.t18 a_6164_n9984.t21 VSS.t31 sky130_fd_pr__res_high_po_0p69 l=12.22
X62 a_n2121_n9699# a_n2577_n10167# VDD.t11 VDD.t10 sky130_fd_pr__pfet_g5v0d10v5 ad=0.2142 pd=1.99 as=0.2142 ps=1.99 w=0.42 l=1
X63 x5.V2.t51 x4.V2.t52 VSS.t44 sky130_fd_pr__res_high_po_0p69 l=12.22
X64 VDD.t165 a_n1825_12142# D03v3.t1 VDD.t96 sky130_fd_pr__pfet_g5v0d10v5 ad=0.24375 pd=1.825 as=0.3975 ps=3.53 w=1.5 l=0.5
X65 x6.V1.t48 x9.V2.t35 VSS.t177 sky130_fd_pr__res_high_po_0p69 l=12.22
X66 VOUT.t4 a_11509_n4916# VSS.t99 sky130_fd_pr__res_high_po_0p69 l=12.22
X67 AVOUT1.t2 a_6164_n4916.t2 VSS.t31 sky130_fd_pr__res_high_po_0p69 l=12.22
X68 x5.V2.t81 x4.V2.t82 VSS.t24 sky130_fd_pr__res_high_po_0p69 l=12.22
X69 ia_opamp_0.V2.t28 a_10959_n8604# VSS.t149 sky130_fd_pr__res_high_po_0p69 l=12.22
X70 VOUT.t14 a_10959_n3536# VSS.t149 sky130_fd_pr__res_high_po_0p69 l=12.22
X71 a_n2577_2313# a_n2603_2366# DVSS.t242 DVSS.t237 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X72 VDD.t118 a_10583_764.t4 x8.V2.t34 VDD.t117 sky130_fd_pr__pfet_g5v0d10v5 ad=5.51 pd=38.58 as=2.755 ps=19.29 w=19 l=1
X73 a_204_12823.t4 a_204_12823.t3 VDD.t130 VDD.t129 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=1
X74 a_n2577_12297# a_n2603_12350# DVSS.t201 DVSS.t196 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X75 x6.V1.t85 x9.V2.t61 VSS.t14 sky130_fd_pr__res_high_po_0p69 l=12.22
X76 x5.V2.t73 x4.V2.t74 VSS.t39 sky130_fd_pr__res_high_po_0p69 l=12.22
X77 x5.V2.t48 x4.V2.t49 VSS.t178 sky130_fd_pr__res_high_po_0p69 l=12.22
X78 DVDD.t7 a_n2559_8407# a_n2603_7358# DVDD.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.12 as=0.2478 ps=2.27 w=0.84 l=0.15
X79 x3.R1.t39 x8.V2.t38 VSS.t150 sky130_fd_pr__res_high_po_0p69 l=12.22
X80 DVSS.t266 a_n2559_919# a_n2121_285# DVSS.t265 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.3975 ps=3.53 w=1.5 l=0.5
X81 a_n2121_n7203# a_n2577_n7671# VDD.t93 VDD.t92 sky130_fd_pr__pfet_g5v0d10v5 ad=0.2142 pd=1.99 as=0.2142 ps=1.99 w=0.42 l=1
X82 a_3720_n9984.t9 D33v3.t4 x5.V2.t58 VSS.t194 sky130_fd_pr__nfet_g5v0d10v5 ad=1.2702 pd=9.34 as=0.6351 ps=4.67 w=4.38 l=1
X83 a_9789_764.t4 a_9789_764.t3 VDD.t30 VDD.t29 sky130_fd_pr__pfet_g5v0d10v5 ad=2.175 pd=15.29 as=4.35 ps=30.58 w=15 l=1
X84 ia_opamp_0.ibias.t1 ia_opamp_0.ibias.t0 VSS.t74 VSS.t73 sky130_fd_pr__nfet_g5v0d10v5 ad=4.4776 pd=31.46 as=4.4776 ps=31.46 w=15.44 l=1
X85 DVSS.t151 a_n2603_9854# a_n2577_9801# DVSS.t146 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X86 a_3720_n4916.t8 D33v3.t5 x4.V2.t61 VSS.t194 sky130_fd_pr__nfet_g5v0d10v5 ad=1.2702 pd=9.34 as=0.6351 ps=4.67 w=4.38 l=1
X87 x3.R1.t82 x8.V2.t59 VSS.t100 sky130_fd_pr__res_high_po_0p69 l=12.22
X88 a_n2121_n7203# a_n2559_n6569# DVSS.t105 DVSS.t104 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X89 VDD.t7 a_16157_764.t2 a_16157_764.t3 VDD.t6 sky130_fd_pr__pfet_g5v0d10v5 ad=4.35 pd=30.58 as=2.175 ps=15.29 w=15 l=1
X90 VDD.t16 a_9789_764.t5 a_10583_764.t0 VDD.t15 sky130_fd_pr__pfet_g5v0d10v5 ad=4.35 pd=30.58 as=2.175 ps=15.29 w=15 l=1
X91 a_n1825_2158# a_n2121_2781# VDD.t181 VDD.t113 sky130_fd_pr__pfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.24375 ps=1.825 w=1.5 l=0.5
X92 DVSS.t256 a_n2559_n4073# a_n2603_n5122# DVSS.t255 sky130_fd_pr__nfet_01v8 ad=0.1176 pd=1.12 as=0.2478 ps=2.27 w=0.84 l=0.15
X93 a_n2559_5911# D3.t0 DVSS.t70 DVSS.t69 sky130_fd_pr__nfet_01v8 ad=0.2478 pd=2.27 as=0.1176 ps=1.12 w=0.84 l=0.15
X94 a_n2559_919# D5.t0 DVSS.t34 DVSS.t33 sky130_fd_pr__nfet_01v8 ad=0.2478 pd=2.27 as=0.1176 ps=1.12 w=0.84 l=0.15
X95 AVOUT2.t19 a_862_n8604# VSS.t122 sky130_fd_pr__res_high_po_0p69 l=12.22
X96 DVSS.t304 VDD.t234 DVSS.t303 DVSS.t302 sky130_fd_pr__nfet_g5v0d10v5 ad=0.19875 pd=2.03 as=0 ps=0 w=0.75 l=1
X97 a_n2121_10269# a_n2559_10903# DVSS.t18 DVSS.t17 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X98 AVOUT1.t30 a_862_n3536# VSS.t122 sky130_fd_pr__res_high_po_0p69 l=12.22
X99 x6.V1.t49 x9.V2.t36 VSS.t150 sky130_fd_pr__res_high_po_0p69 l=12.22
X100 VDD.t159 DVSS.t308 VDD.t158 VDD.t157 sky130_fd_pr__pfet_g5v0d10v5 ad=0.265 pd=2.53 as=0 ps=0 w=1 l=1
X101 DVSS.t200 a_n2603_12350# a_n2577_12297# DVSS.t196 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X102 a_16157_764.t1 a_16157_764.t0 VDD.t5 VDD.t4 sky130_fd_pr__pfet_g5v0d10v5 ad=2.175 pd=15.29 as=4.35 ps=30.58 w=15 l=1
X103 AVOUT2.t34 a_3720_n9984.t14 VSS.t32 sky130_fd_pr__res_high_po_0p69 l=12.22
X104 x6.V1.t25 x9.V2.t13 VSS.t100 sky130_fd_pr__res_high_po_0p69 l=12.22
X105 DVDD.t23 a_n2559_n6569# a_n2603_n7618# DVDD.t22 sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.12 as=0.2478 ps=2.27 w=0.84 l=0.15
X106 a_n2121_n9699# a_n2559_n9065# DVSS.t167 DVSS.t166 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X107 x5.V2.t16 D33v3.t6 a_3720_n9984.t8 VSS.t86 sky130_fd_pr__nfet_g5v0d10v5 ad=0.6351 pd=4.67 as=0.6351 ps=4.67 w=4.38 l=1
X108 AVOUT1.t3 a_3720_n4916.t0 VSS.t32 sky130_fd_pr__res_high_po_0p69 l=12.22
X109 DVSS.t165 a_n2559_n9065# a_n2121_n9699# DVSS.t164 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X110 x3.R1.t22 x8.V2.t18 VSS.t116 sky130_fd_pr__res_high_po_0p69 l=12.22
X111 DVSS.t191 a_n1825_12142# D03v3.t0 DVSS.t190 sky130_fd_pr__nfet_g5v0d10v5 ad=0.121875 pd=1.075 as=0.19875 ps=2.03 w=0.75 l=0.5
X112 a_6164_n9984.t15 D43v3.t6 x5.V2.t83 VSS.t244 sky130_fd_pr__nfet_g5v0d10v5 ad=0.638 pd=4.69 as=0.638 ps=4.69 w=4.4 l=1
X113 x4.V2.t17 D33v3.t7 a_3720_n4916.t7 VSS.t86 sky130_fd_pr__nfet_g5v0d10v5 ad=0.6351 pd=4.67 as=0.6351 ps=4.67 w=4.38 l=1
X114 a_n2559_3415# D4.t0 DVSS.t49 DVSS.t48 sky130_fd_pr__nfet_01v8 ad=0.2478 pd=2.27 as=0.1176 ps=1.12 w=0.84 l=0.15
X115 DVSS.t301 VDD.t235 DVSS.t300 DVSS.t299 sky130_fd_pr__nfet_g5v0d10v5 ad=0.19875 pd=2.03 as=0 ps=0 w=0.75 l=1
X116 x3.R1.t41 x8.V2.t40 VSS.t63 sky130_fd_pr__res_high_po_0p69 l=12.22
X117 ia_opamp_0.V2.t2 a_16261_n9984.t2 VSS.t33 sky130_fd_pr__res_high_po_0p69 l=12.22
X118 a_n2121_12765# a_n2559_13399# DVSS.t226 DVSS.t225 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X119 x5.V2.t17 D33v3.t8 a_3720_n9984.t7 VSS.t87 sky130_fd_pr__nfet_g5v0d10v5 ad=0.6351 pd=4.67 as=0.6351 ps=4.67 w=4.38 l=1
X120 a_6164_n4916.t16 D43v3.t7 x4.V2.t85 VSS.t244 sky130_fd_pr__nfet_g5v0d10v5 ad=0.638 pd=4.69 as=0.638 ps=4.69 w=4.4 l=1
X121 x5.V2.t11 x4.V2.t12 VSS.t60 sky130_fd_pr__res_high_po_0p69 l=12.22
X122 x4.V2.t42 D33v3.t9 a_3720_n4916.t6 VSS.t87 sky130_fd_pr__nfet_g5v0d10v5 ad=0.6351 pd=4.67 as=0.6351 ps=4.67 w=4.38 l=1
X123 VOUT.t27 a_16261_n4916.t13 VSS.t33 sky130_fd_pr__res_high_po_0p69 l=12.22
X124 a_n2577_4809# a_n2603_4862# DVSS.t181 DVSS.t176 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X125 x5.V2.t31 x4.V2.t30 VSS.t63 sky130_fd_pr__res_high_po_0p69 l=12.22
X126 a_n2577_14793# a_n2603_14846# DVSS.t175 DVSS.t170 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X127 x3.R1.t11 x8.V2.t10 VSS.t61 sky130_fd_pr__res_high_po_0p69 l=12.22
X128 amp_biases_0.ibias1.t1 amp_biases_0.ibias1.t0 VSS.t50 VSS.t49 sky130_fd_pr__nfet_g5v0d10v5 ad=4.4776 pd=31.46 as=4.4776 ps=31.46 w=15.44 l=1
X129 x3.R1.t12 x8.V2.t11 VSS.t62 sky130_fd_pr__res_high_po_0p69 l=12.22
X130 x6.V1.t28 x9.V2.t15 VSS.t116 sky130_fd_pr__res_high_po_0p69 l=12.22
X131 x5.V2.t29 x4.V2.t28 VSS.t112 sky130_fd_pr__res_high_po_0p69 l=12.22
X132 a_16261_n9984.t26 D93v3.t4 x6.V1.t61 VSS.t202 sky130_fd_pr__nfet_g5v0d10v5 ad=0.638 pd=4.69 as=0.638 ps=4.69 w=4.4 l=1
X133 AVOUT2.t0 a_6164_n9984.t0 VSS.t3 sky130_fd_pr__res_high_po_0p69 l=12.22
X134 a_10047_764.t0 x8.V2.t70 a_9789_764.t0 VSS.t201 sky130_fd_pr__nfet_g5v0d10v5 ad=4.785 pd=33.58 as=4.785 ps=33.58 w=16.5 l=1
X135 a_4215_764.t3 a_3421_764.t5 VDD.t122 VDD.t121 sky130_fd_pr__pfet_g5v0d10v5 ad=2.175 pd=15.29 as=4.35 ps=30.58 w=15 l=1
X136 x5.V2.t46 x4.V2.t48 VSS.t152 sky130_fd_pr__res_high_po_0p69 l=12.22
X137 x6.V1.t16 x9.V2.t8 VSS.t63 sky130_fd_pr__res_high_po_0p69 l=12.22
X138 a_16261_n4916.t26 D93v3.t5 x3.R1.t78 VSS.t202 sky130_fd_pr__nfet_g5v0d10v5 ad=0.638 pd=4.69 as=0.638 ps=4.69 w=4.4 l=1
X139 AVOUT1.t17 a_6164_n4916.t19 VSS.t3 sky130_fd_pr__res_high_po_0p69 l=12.22
X140 DVSS.t125 a_n2559_15895# a_n2121_15261# DVSS.t124 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.3975 ps=3.53 w=1.5 l=0.5
X141 DVSS.t298 VDD.t236 DVSS.t297 DVSS.t296 sky130_fd_pr__nfet_g5v0d10v5 ad=0.19875 pd=2.03 as=0 ps=0 w=0.75 l=1
X142 AVOUT2.t33 a_6164_n9984.t28 VSS.t34 sky130_fd_pr__res_high_po_0p69 l=12.22
X143 a_495_764.t2 ia_opamp_0.V2.t38 a_237_764.t4 VSS.t115 sky130_fd_pr__nfet_g5v0d10v5 ad=4.785 pd=33.58 as=4.785 ps=33.58 w=16.5 l=1
X144 VDD.t69 a_3421_764.t3 a_3421_764.t4 VDD.t68 sky130_fd_pr__pfet_g5v0d10v5 ad=4.35 pd=30.58 as=2.175 ps=15.29 w=15 l=1
X145 DVSS.t234 a_n2603_7358# a_n2577_7305# DVSS.t229 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.3975 ps=3.53 w=1.5 l=0.5
X146 AVOUT1.t4 a_6164_n4916.t3 VSS.t34 sky130_fd_pr__res_high_po_0p69 l=12.22
X147 a_3720_n9984.t6 D33v3.t10 x5.V2.t41 VSS.t159 sky130_fd_pr__nfet_g5v0d10v5 ad=0.6351 pd=4.67 as=0.6351 ps=4.67 w=4.38 l=1
X148 VDD.t144 a_7399_764.t4 AVOUT2.t23 VDD.t143 sky130_fd_pr__pfet_g5v0d10v5 ad=5.51 pd=38.58 as=2.755 ps=19.29 w=19 l=1
X149 a_n2559_8407# D2.t0 DVSS.t55 DVSS.t54 sky130_fd_pr__nfet_01v8 ad=0.2478 pd=2.27 as=0.1176 ps=1.12 w=0.84 l=0.15
X150 x6.V1.t62 x9.V2.t43 VSS.t61 sky130_fd_pr__res_high_po_0p69 l=12.22
X151 x5.V2.t32 x4.V2.t31 VSS.t118 sky130_fd_pr__res_high_po_0p69 l=12.22
X152 a_3720_n4916.t5 D33v3.t11 x4.V2.t43 VSS.t159 sky130_fd_pr__nfet_g5v0d10v5 ad=0.6351 pd=4.67 as=0.6351 ps=4.67 w=4.38 l=1
X153 a_4215_764.t0 V2.t0 a_3679_764.t2 VSS.t84 sky130_fd_pr__nfet_g5v0d10v5 ad=4.785 pd=33.58 as=4.785 ps=33.58 w=16.5 l=1
X154 x5.V2.t87 x4.V2.t88 VSS.t170 sky130_fd_pr__res_high_po_0p69 l=12.22
X155 DVSS.t3 a_n1825_n10322# D93v3.t0 DVSS.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=0.121875 pd=1.075 as=0.19875 ps=2.03 w=0.75 l=0.5
X156 x5.V2.t42 x4.V2.t44 VSS.t142 sky130_fd_pr__res_high_po_0p69 l=12.22
X157 x6.V1.t42 x9.V2.t29 VSS.t62 sky130_fd_pr__res_high_po_0p69 l=12.22
X158 x3.R1.t19 x8.V2.t15 VSS.t91 sky130_fd_pr__res_high_po_0p69 l=12.22
X159 ia_opamp_0.V2.t4 a_16261_n9984.t4 VSS.t56 sky130_fd_pr__res_high_po_0p69 l=12.22
X160 a_3421_764.t2 a_3421_764.t1 VDD.t91 VDD.t90 sky130_fd_pr__pfet_g5v0d10v5 ad=2.175 pd=15.29 as=4.35 ps=30.58 w=15 l=1
X161 VOUT.t2 a_16261_n4916.t0 VSS.t56 sky130_fd_pr__res_high_po_0p69 l=12.22
X162 DVSS.t5 a_n1825_n338# D53v3.t0 DVSS.t4 sky130_fd_pr__nfet_g5v0d10v5 ad=0.121875 pd=1.075 as=0.19875 ps=2.03 w=0.75 l=0.5
X163 a_1031_764.t1 G.t0 a_495_764.t0 VSS.t122 sky130_fd_pr__nfet_g5v0d10v5 ad=4.785 pd=33.58 as=4.785 ps=33.58 w=16.5 l=1
X164 DVSS.t150 a_n2603_9854# a_n2577_9801# DVSS.t146 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.3975 ps=3.53 w=1.5 l=0.5
X165 DVSS.t29 a_n1825_9646# D13v3.t0 DVSS.t28 sky130_fd_pr__nfet_g5v0d10v5 ad=0.121875 pd=1.075 as=0.19875 ps=2.03 w=0.75 l=0.5
X166 DVSS.t143 a_n2603_n2626# a_n2577_n2679# DVSS.t138 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X167 DVDD.t31 a_n2559_n9065# a_n2603_n10114# DVDD.t30 sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.12 as=0.2478 ps=2.27 w=0.84 l=0.15
X168 ia_opamp_0.V2.t16 a_13817_n9984.t1 VSS.t161 sky130_fd_pr__res_high_po_0p69 l=12.22
X169 x5.V2.t74 x4.V2.t75 VSS.t35 sky130_fd_pr__res_high_po_0p69 l=12.22
X170 x3.R1.t34 x8.V2.t29 VSS.t142 sky130_fd_pr__res_high_po_0p69 l=12.22
X171 VDD.t112 a_9789_764.t1 a_9789_764.t2 VDD.t111 sky130_fd_pr__pfet_g5v0d10v5 ad=4.35 pd=30.58 as=2.175 ps=15.29 w=15 l=1
X172 a_n2121_285# a_n2559_919# DVSS.t264 DVSS.t263 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X173 x3.R1.t14 x8.V2.t13 VSS.t44 sky130_fd_pr__res_high_po_0p69 l=12.22
X174 VOUT.t17 a_13817_n4916.t4 VSS.t161 sky130_fd_pr__res_high_po_0p69 l=12.22
X175 DVSS.t66 a_n2559_5911# a_n2121_5277# DVSS.t65 sky130_fd_pr__nfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.21 ps=1.78 w=1.5 l=0.5
X176 x3.R1.t81 x8.V2.t58 VSS.t143 sky130_fd_pr__res_high_po_0p69 l=12.22
X177 VDD.t61 a_6605_764.t5 a_7399_764.t1 VDD.t60 sky130_fd_pr__pfet_g5v0d10v5 ad=4.35 pd=30.58 as=2.175 ps=15.29 w=15 l=1
X178 VDD.t132 a_204_12823.t5 amp_biases_0.ibias1.t3 VDD.t131 sky130_fd_pr__pfet_g5v0d10v5 ad=2.175 pd=15.29 as=2.175 ps=15.29 w=15 l=1
X179 a_n2577_9801# a_n2121_10269# VDD.t128 VDD.t127 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1365 pd=1.49 as=0.1113 ps=1.37 w=0.42 l=1
X180 DVSS.t202 D7.t0 sky130_fd_pr__diode_pw2nd_11v0 perim=3.16e+06 area=6.072e+11
X181 x6.V1.t88 x9.V2.t64 VSS.t91 sky130_fd_pr__res_high_po_0p69 l=12.22
X182 VDD.t162 DVSS.t309 VDD.t161 VDD.t160 sky130_fd_pr__pfet_g5v0d10v5 ad=0.265 pd=2.53 as=0 ps=0 w=1 l=1
X183 a_n2559_n9065# D9.t1 DVSS.t169 DVSS.t168 sky130_fd_pr__nfet_01v8 ad=0.2478 pd=2.27 as=0.1176 ps=1.12 w=0.84 l=0.15
X184 a_16150_281.t0 VOUT.t29 VSS.t228 sky130_fd_pr__res_high_po_0p69 l=3.2
X185 VDD.t138 a_204_12823.t6 amp_biases_0.ibias5.t3 VDD.t137 sky130_fd_pr__pfet_g5v0d10v5 ad=4.35 pd=30.58 as=2.175 ps=15.29 w=15 l=1
X186 x5.V2.t25 D23v3.t2 a_2308_n9984.t3 VSS.t123 sky130_fd_pr__nfet_g5v0d10v5 ad=0.67425 pd=4.94 as=1.3485 ps=9.88 w=4.65 l=1
X187 a_n1825_n2834# a_n2121_n2211# VDD.t89 VDD.t88 sky130_fd_pr__pfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.24375 ps=1.825 w=1.5 l=0.5
X188 x4.V2.t35 D23v3.t3 a_2308_n4916.t3 VSS.t123 sky130_fd_pr__nfet_g5v0d10v5 ad=0.67425 pd=4.94 as=1.3485 ps=9.88 w=4.65 l=1
X189 AVOUT2.t10 a_6164_n9984.t3 VSS.t105 sky130_fd_pr__res_high_po_0p69 l=12.22
X190 amp_biases_0.ibias2.t1 amp_biases_0.ibias2.t0 VSS.t219 VSS.t218 sky130_fd_pr__nfet_g5v0d10v5 ad=4.4776 pd=31.46 as=4.4776 ps=31.46 w=15.44 l=1
X191 a_n2577_n10167# a_n2603_n10114# DVSS.t26 DVSS.t22 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X192 a_n2577_n183# a_n2603_n130# DVSS.t187 DVSS.t182 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X193 x6.V1.t32 x9.V2.t19 VSS.t142 sky130_fd_pr__res_high_po_0p69 l=12.22
X194 AVOUT1.t28 a_6164_n4916.t25 VSS.t105 sky130_fd_pr__res_high_po_0p69 l=12.22
X195 DVSS.t45 a_n2559_8407# a_n2121_7773# DVSS.t44 sky130_fd_pr__nfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.21 ps=1.78 w=1.5 l=0.5
X196 DVSS.t212 a_n2559_3415# a_n2121_2781# DVSS.t211 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.3975 ps=3.53 w=1.5 l=0.5
X197 x6.V1.t33 x9.V2.t20 VSS.t143 sky130_fd_pr__res_high_po_0p69 l=12.22
X198 x6.V1.t11 x9.V2.t5 VSS.t44 sky130_fd_pr__res_high_po_0p69 l=12.22
X199 AVOUT2.t1 a_3720_n9984.t0 VSS.t37 sky130_fd_pr__res_high_po_0p69 l=12.22
X200 a_7399_764.t0 a_6605_764.t6 VDD.t183 VDD.t182 sky130_fd_pr__pfet_g5v0d10v5 ad=2.175 pd=15.29 as=4.35 ps=30.58 w=15 l=1
X201 VDD.t48 a_6605_764.t0 a_6605_764.t1 VDD.t47 sky130_fd_pr__pfet_g5v0d10v5 ad=4.35 pd=30.58 as=2.175 ps=15.29 w=15 l=1
X202 a_n2577_12297# a_n2121_12765# VDD.t99 VDD.t98 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1365 pd=1.49 as=0.1113 ps=1.37 w=0.42 l=1
X203 ia_opamp_0.V2.t14 a_16261_n9984.t9 VSS.t113 sky130_fd_pr__res_high_po_0p69 l=12.22
X204 AVOUT1.t24 a_3720_n4916.t14 VSS.t37 sky130_fd_pr__res_high_po_0p69 l=12.22
X205 a_3414_281.t0 AVOUT1.t11 VSS.t93 sky130_fd_pr__res_high_po_0p69 l=3.2
X206 VDD.t204 DVSS.t310 VDD.t203 VDD.t202 sky130_fd_pr__pfet_g5v0d10v5 ad=0.265 pd=2.53 as=0 ps=0 w=1 l=1
X207 x3.R1.t9 x8.V2.t8 VSS.t57 sky130_fd_pr__res_high_po_0p69 l=12.22
X208 a_n2559_10903# D1.t0 DVSS.t1 DVSS.t0 sky130_fd_pr__nfet_01v8 ad=0.2478 pd=2.27 as=0.1176 ps=1.12 w=0.84 l=0.15
X209 a_n2121_5277# a_n2577_4809# VDD.t199 VDD.t198 sky130_fd_pr__pfet_g5v0d10v5 ad=0.2142 pd=1.99 as=0.2142 ps=1.99 w=0.42 l=1
X210 VOUT.t9 a_16261_n4916.t3 VSS.t113 sky130_fd_pr__res_high_po_0p69 l=12.22
X211 VDD.t136 a_12973_764.t5 a_13767_764.t1 VDD.t135 sky130_fd_pr__pfet_g5v0d10v5 ad=4.35 pd=30.58 as=2.175 ps=15.29 w=15 l=1
X212 a_1412_n9984# D13v3.t2 x5.V2.t91 VSS.t154 sky130_fd_pr__nfet_g5v0d10v5 ad=1.4123 pd=10.32 as=0.70615 ps=5.16 w=4.87 l=1
X213 amp_biases_0.ibias1.t2 a_204_12823.t7 VDD.t140 VDD.t139 sky130_fd_pr__pfet_g5v0d10v5 ad=2.175 pd=15.29 as=2.175 ps=15.29 w=15 l=1
X214 a_1412_n4916# D13v3.t3 x4.V2.t40 VSS.t154 sky130_fd_pr__nfet_g5v0d10v5 ad=1.4123 pd=10.32 as=0.70615 ps=5.16 w=4.87 l=1
X215 DVSS.t64 a_n2559_5911# a_n2121_5277# DVSS.t63 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.3975 ps=3.53 w=1.5 l=0.5
X216 x5.V2.t71 x4.V2.t72 VSS.t79 sky130_fd_pr__res_high_po_0p69 l=12.22
X217 a_6863_764.t2 x5.V2.t94 a_6605_764.t4 VSS.t129 sky130_fd_pr__nfet_g5v0d10v5 ad=4.785 pd=33.58 as=4.785 ps=33.58 w=16.5 l=1
X218 x5.V2.t44 x4.V2.t46 VSS.t114 sky130_fd_pr__res_high_po_0p69 l=12.22
X219 DVDD.t35 a_n2559_3415# a_n2603_2366# DVDD.t34 sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.12 as=0.2478 ps=2.27 w=0.84 l=0.15
X220 x6.V1.t44 x9.V2.t31 VSS.t57 sky130_fd_pr__res_high_po_0p69 l=12.22
X221 AVOUT2.t30 a_1412_n9984# VSS.t241 sky130_fd_pr__res_high_po_0p69 l=12.22
X222 a_n2121_7773# a_n2577_7305# VDD.t191 VDD.t190 sky130_fd_pr__pfet_g5v0d10v5 ad=0.2142 pd=1.99 as=0.2142 ps=1.99 w=0.42 l=1
X223 a_n2121_n2211# a_n2577_n2679# VDD.t81 VDD.t80 sky130_fd_pr__pfet_g5v0d10v5 ad=0.2142 pd=1.99 as=0.2142 ps=1.99 w=0.42 l=1
X224 AVOUT1.t37 a_1412_n4916# VSS.t241 sky130_fd_pr__res_high_po_0p69 l=12.22
X225 VDD.t59 a_12973_764.t0 a_12973_764.t1 VDD.t58 sky130_fd_pr__pfet_g5v0d10v5 ad=4.35 pd=30.58 as=2.175 ps=15.29 w=15 l=1
X226 DVSS.t186 a_n2603_n130# a_n2577_n183# DVSS.t182 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X227 x5.V2.t84 D43v3.t8 a_6164_n9984.t14 VSS.t47 sky130_fd_pr__nfet_g5v0d10v5 ad=0.638 pd=4.69 as=0.638 ps=4.69 w=4.4 l=1
X228 x8.V2.t35 a_10583_764.t5 VDD.t120 VDD.t119 sky130_fd_pr__pfet_g5v0d10v5 ad=2.755 pd=19.29 as=5.51 ps=38.58 w=19 l=1
X229 a_n2121_n2211# a_n2559_n1577# DVSS.t83 DVSS.t82 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X230 VDD.t142 a_204_12823.t8 ia_opamp_0.ibias.t3 VDD.t141 sky130_fd_pr__pfet_g5v0d10v5 ad=2.175 pd=15.29 as=2.175 ps=15.29 w=15 l=1
X231 x5.V2.t56 x4.V2.t57 VSS.t116 sky130_fd_pr__res_high_po_0p69 l=12.22
X232 AVOUT2.t25 a_6164_n9984.t23 VSS.t208 sky130_fd_pr__res_high_po_0p69 l=12.22
X233 x5.V2.t14 x4.V2.t15 VSS.t61 sky130_fd_pr__res_high_po_0p69 l=12.22
X234 x5.V2.t69 x4.V2.t70 VSS.t8 sky130_fd_pr__res_high_po_0p69 l=12.22
X235 x4.V2.t9 D43v3.t9 a_6164_n4916.t15 VSS.t47 sky130_fd_pr__nfet_g5v0d10v5 ad=0.638 pd=4.69 as=0.638 ps=4.69 w=4.4 l=1
X236 x3.R1.t87 x8.V2.t64 VSS.t174 sky130_fd_pr__res_high_po_0p69 l=12.22
X237 AVOUT1.t35 a_6164_n4916.t29 VSS.t208 sky130_fd_pr__res_high_po_0p69 l=12.22
X238 ia_opamp_0.V2.t8 a_16261_n9984.t7 VSS.t92 sky130_fd_pr__res_high_po_0p69 l=12.22
X239 x5.V2.t8 D43v3.t10 a_6164_n9984.t13 VSS.t48 sky130_fd_pr__nfet_g5v0d10v5 ad=0.638 pd=4.69 as=0.638 ps=4.69 w=4.4 l=1
X240 a_12405_n9984.t4 D73v3.t4 x6.V1.t17 VSS.t76 sky130_fd_pr__nfet_g5v0d10v5 ad=0.67425 pd=4.94 as=0.67425 ps=4.94 w=4.65 l=1
X241 a_n2121_7773# a_n2559_8407# DVSS.t47 DVSS.t46 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X242 DVDD.t13 a_n2559_5911# a_n2603_4862# DVDD.t12 sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.12 as=0.2478 ps=2.27 w=0.84 l=0.15
X243 a_n1825_n2834# a_n2121_n2211# DVSS.t75 DVSS.t74 sky130_fd_pr__nfet_g5v0d10v5 ad=0.19875 pd=2.03 as=0.121875 ps=1.075 w=0.75 l=0.5
X244 DVSS.t43 a_n2559_8407# a_n2603_7358# DVSS.t42 sky130_fd_pr__nfet_01v8 ad=0.1176 pd=1.12 as=0.2478 ps=2.27 w=0.84 l=0.15
X245 a_n1825_n5330# a_n2121_n4707# VDD.t225 VDD.t188 sky130_fd_pr__pfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.24375 ps=1.825 w=1.5 l=0.5
X246 a_12405_n4916.t5 D73v3.t5 x3.R1.t16 VSS.t76 sky130_fd_pr__nfet_g5v0d10v5 ad=0.67425 pd=4.94 as=0.67425 ps=4.94 w=4.65 l=1
X247 x4.V2.t10 D43v3.t11 a_6164_n4916.t14 VSS.t48 sky130_fd_pr__nfet_g5v0d10v5 ad=0.638 pd=4.69 as=0.638 ps=4.69 w=4.4 l=1
X248 DVSS.t108 D1.t1 sky130_fd_pr__diode_pw2nd_11v0 perim=3.16e+06 area=6.072e+11
X249 VOUT.t3 a_16261_n4916.t1 VSS.t92 sky130_fd_pr__res_high_po_0p69 l=12.22
X250 x5.V2.t55 x4.V2.t56 VSS.t132 sky130_fd_pr__res_high_po_0p69 l=12.22
X251 x5.V2.t1 x4.V2.t1 VSS.t4 sky130_fd_pr__res_high_po_0p69 l=12.22
X252 ia_opamp_0.ibias.t2 a_204_12823.t9 VDD.t36 VDD.t35 sky130_fd_pr__pfet_g5v0d10v5 ad=2.175 pd=15.29 as=4.35 ps=30.58 w=15 l=1
X253 ia_opamp_0.V2.t19 a_13817_n9984.t3 VSS.t117 sky130_fd_pr__res_high_po_0p69 l=12.22
X254 a_6598_281.t1 a_7399_764.t2 sky130_fd_pr__cap_mim_m3_1 l=6.9 w=6.9
X255 x5.V2.t93 x4.V2.t93 VSS.t7 sky130_fd_pr__res_high_po_0p69 l=12.22
X256 x3.R1.t84 x8.V2.t61 VSS.t141 sky130_fd_pr__res_high_po_0p69 l=12.22
X257 DVSS.t295 VDD.t237 DVSS.t294 DVSS.t293 sky130_fd_pr__nfet_g5v0d10v5 ad=0.19875 pd=2.03 as=0 ps=0 w=0.75 l=1
X258 DVDD.t19 a_n2559_n1577# a_n2603_n2626# DVDD.t18 sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.12 as=0.2478 ps=2.27 w=0.84 l=0.15
X259 a_n2121_n4707# a_n2559_n4073# DVSS.t254 DVSS.t253 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X260 VOUT.t10 a_13817_n4916.t1 VSS.t117 sky130_fd_pr__res_high_po_0p69 l=12.22
X261 x3.R1.t6 x8.V2.t6 VSS.t43 sky130_fd_pr__res_high_po_0p69 l=12.22
X262 ia_opamp_0.V2.t17 a_16261_n9984.t10 VSS.t156 sky130_fd_pr__res_high_po_0p69 l=12.22
X263 DVSS.t252 a_n2559_n4073# a_n2121_n4707# DVSS.t251 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X264 x3.R1.t52 x8.V2.t52 VSS.t217 sky130_fd_pr__res_high_po_0p69 l=12.22
X265 x6.V1.t46 x9.V2.t33 VSS.t174 sky130_fd_pr__res_high_po_0p69 l=12.22
X266 VOUT.t15 a_16261_n4916.t5 VSS.t156 sky130_fd_pr__res_high_po_0p69 l=12.22
X267 a_n2559_13399# D0.t0 DVSS.t136 DVSS.t135 sky130_fd_pr__nfet_01v8 ad=0.2478 pd=2.27 as=0.1176 ps=1.12 w=0.84 l=0.15
X268 VDD.t9 a_n1825_n338# D53v3.t1 VDD.t8 sky130_fd_pr__pfet_g5v0d10v5 ad=0.24375 pd=1.825 as=0.3975 ps=3.53 w=1.5 l=0.5
X269 x6.V1.t70 D93v3.t6 a_16261_n9984.t25 VSS.t227 sky130_fd_pr__nfet_g5v0d10v5 ad=0.638 pd=4.69 as=0.638 ps=4.69 w=4.4 l=1
X270 VDD.t44 a_16157_764.t6 a_16951_764.t2 VDD.t43 sky130_fd_pr__pfet_g5v0d10v5 ad=4.35 pd=30.58 as=2.175 ps=15.29 w=15 l=1
X271 VDD.t164 a_237_764.t5 a_1031_764.t3 VDD.t163 sky130_fd_pr__pfet_g5v0d10v5 ad=4.35 pd=30.58 as=2.175 ps=15.29 w=15 l=1
X272 VDD.t32 a_n1825_9646# D13v3.t1 VDD.t31 sky130_fd_pr__pfet_g5v0d10v5 ad=0.24375 pd=1.825 as=0.3975 ps=3.53 w=1.5 l=0.5
X273 DVSS.t292 VDD.t238 DVSS.t291 DVSS.t290 sky130_fd_pr__nfet_g5v0d10v5 ad=0.19875 pd=2.03 as=0 ps=0 w=0.75 l=1
X274 a_n1825_n7826# a_n2121_n7203# VDD.t125 VDD.t84 sky130_fd_pr__pfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.24375 ps=1.825 w=1.5 l=0.5
X275 a_n1825_n10322# a_n2121_n9699# VDD.t14 VDD.t0 sky130_fd_pr__pfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.24375 ps=1.825 w=1.5 l=0.5
X276 x3.R1.t77 D93v3.t7 a_16261_n4916.t22 VSS.t227 sky130_fd_pr__nfet_g5v0d10v5 ad=0.638 pd=4.69 as=0.638 ps=4.69 w=4.4 l=1
X277 x5.V2.t30 x4.V2.t29 VSS.t137 sky130_fd_pr__res_high_po_0p69 l=12.22
X278 DVSS.t224 a_n2559_13399# a_n2121_12765# DVSS.t223 sky130_fd_pr__nfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.21 ps=1.78 w=1.5 l=0.5
X279 ibias.t0 sky130_fd_sc_hvl__lsbuflv2hv_1_0[10].X.t2 a_2622_12748.t0 VSS.t235 sky130_fd_pr__nfet_g5v0d10v5 ad=4.4776 pd=31.46 as=2.2388 ps=15.73 w=15.44 l=1
X280 a_12966_281.t1 a_13767_764.t2 sky130_fd_pr__cap_mim_m3_1 l=6.9 w=6.9
X281 AVOUT2.t9 a_6164_n9984.t2 VSS.t103 sky130_fd_pr__res_high_po_0p69 l=12.22
X282 DVSS.t180 a_n2603_4862# a_n2577_4809# DVSS.t176 sky130_fd_pr__nfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.21 ps=1.78 w=1.5 l=0.5
X283 a_6164_n9984.t12 D43v3.t12 x5.V2.t61 VSS.t196 sky130_fd_pr__nfet_g5v0d10v5 ad=0.638 pd=4.69 as=0.638 ps=4.69 w=4.4 l=1
X284 a_n2577_9801# a_n2603_9854# DVSS.t149 DVSS.t146 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X285 x6.V1.t31 x9.V2.t18 VSS.t141 sky130_fd_pr__res_high_po_0p69 l=12.22
X286 AVOUT1.t21 a_6164_n4916.t21 VSS.t103 sky130_fd_pr__res_high_po_0p69 l=12.22
X287 DVSS.t41 a_n2559_8407# a_n2121_7773# DVSS.t40 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.3975 ps=3.53 w=1.5 l=0.5
X288 a_6164_n4916.t13 D43v3.t13 x4.V2.t63 VSS.t196 sky130_fd_pr__nfet_g5v0d10v5 ad=0.638 pd=4.69 as=0.638 ps=4.69 w=4.4 l=1
X289 a_1031_764.t0 a_237_764.t6 VDD.t18 VDD.t17 sky130_fd_pr__pfet_g5v0d10v5 ad=2.175 pd=15.29 as=4.35 ps=30.58 w=15 l=1
X290 DVSS.t103 a_n2559_n6569# a_n2121_n7203# DVSS.t102 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X291 x6.V1.t34 x9.V2.t21 VSS.t43 sky130_fd_pr__res_high_po_0p69 l=12.22
X292 x6.V1.t65 x9.V2.t47 VSS.t217 sky130_fd_pr__res_high_po_0p69 l=12.22
X293 a_6164_n9984.t11 D43v3.t14 x5.V2.t62 VSS.t197 sky130_fd_pr__nfet_g5v0d10v5 ad=0.638 pd=4.69 as=0.638 ps=4.69 w=4.4 l=1
X294 DVSS.t269 ena.t0 sky130_fd_pr__diode_pw2nd_11v0 perim=3.16e+06 area=6.072e+11
X295 a_9782_281.t1 a_10583_764.t2 sky130_fd_pr__cap_mim_m3_1 l=6.9 w=6.9
X296 x5.V2.t3 x4.V2.t3 VSS.t13 sky130_fd_pr__res_high_po_0p69 l=12.22
X297 a_n2559_15895# ena.t1 DVSS.t271 DVSS.t270 sky130_fd_pr__nfet_01v8 ad=0.2478 pd=2.27 as=0.1176 ps=1.12 w=0.84 l=0.15
X298 a_6164_n4916.t12 D43v3.t15 x4.V2.t83 VSS.t197 sky130_fd_pr__nfet_g5v0d10v5 ad=0.638 pd=4.69 as=0.638 ps=4.69 w=4.4 l=1
X299 AVOUT2.t12 a_6164_n9984.t18 VSS.t138 sky130_fd_pr__res_high_po_0p69 l=12.22
X300 x5.V2.t79 x4.V2.t80 VSS.t64 sky130_fd_pr__res_high_po_0p69 l=12.22
X301 DVSS.t16 a_n2559_10903# a_n2121_10269# DVSS.t15 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.3975 ps=3.53 w=1.5 l=0.5
X302 a_12966_281.t0 x9.V2.t17 VSS.t140 sky130_fd_pr__res_high_po_0p69 l=3.2
X303 x3.R1.t47 x8.V2.t47 VSS.t126 sky130_fd_pr__res_high_po_0p69 l=12.22
X304 AVOUT1.t18 a_6164_n4916.t20 VSS.t138 sky130_fd_pr__res_high_po_0p69 l=12.22
X305 VSS.t68 amp_biases_0.ibias2.t4 a_6863_764.t0 VSS.t67 sky130_fd_pr__nfet_g5v0d10v5 ad=4.4776 pd=31.46 as=4.4776 ps=31.46 w=15.44 l=1
X306 a_n1825_12142# a_n2121_12765# VDD.t97 VDD.t96 sky130_fd_pr__pfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.24375 ps=1.825 w=1.5 l=0.5
X307 DVSS.t289 VDD.t239 DVSS.t288 DVSS.t287 sky130_fd_pr__nfet_g5v0d10v5 ad=0.19875 pd=2.03 as=0 ps=0 w=0.75 l=1
X308 DVSS.t233 a_n2603_7358# a_n2577_7305# DVSS.t229 sky130_fd_pr__nfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.21 ps=1.78 w=1.5 l=0.5
X309 DVSS.t241 a_n2603_2366# a_n2577_2313# DVSS.t237 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.3975 ps=3.53 w=1.5 l=0.5
X310 DVSS.t145 a_n1825_2158# D43v3.t0 DVSS.t144 sky130_fd_pr__nfet_g5v0d10v5 ad=0.121875 pd=1.075 as=0.19875 ps=2.03 w=0.75 l=0.5
X311 DVSS.t286 VDD.t240 DVSS.t285 DVSS.t284 sky130_fd_pr__nfet_g5v0d10v5 ad=0.19875 pd=2.03 as=0 ps=0 w=0.75 l=1
X312 x3.R1.t51 x8.V2.t51 VSS.t184 sky130_fd_pr__res_high_po_0p69 l=12.22
X313 ia_opamp_0.V2.t23 a_16261_n9984.t13 VSS.t179 sky130_fd_pr__res_high_po_0p69 l=12.22
X314 a_16261_n9984.t24 D93v3.t8 x6.V1.t71 VSS.t185 sky130_fd_pr__nfet_g5v0d10v5 ad=0.638 pd=4.69 as=0.638 ps=4.69 w=4.4 l=1
X315 x3.R1.t13 x8.V2.t12 VSS.t64 sky130_fd_pr__res_high_po_0p69 l=12.22
X316 VOUT.t20 a_16261_n4916.t8 VSS.t179 sky130_fd_pr__res_high_po_0p69 l=12.22
X317 a_16261_n4916.t21 D93v3.t9 x3.R1.t76 VSS.t185 sky130_fd_pr__nfet_g5v0d10v5 ad=0.638 pd=4.69 as=0.638 ps=4.69 w=4.4 l=1
X318 x3.R1.t25 x8.V2.t21 VSS.t102 sky130_fd_pr__res_high_po_0p69 l=12.22
X319 x5.V2.t43 x4.V2.t45 VSS.t164 sky130_fd_pr__res_high_po_0p69 l=12.22
X320 a_n1825_n5330# a_n2121_n4707# DVSS.t306 DVSS.t305 sky130_fd_pr__nfet_g5v0d10v5 ad=0.19875 pd=2.03 as=0.121875 ps=1.075 w=0.75 l=0.5
X321 a_16261_n9984.t23 D93v3.t10 x6.V1.t55 VSS.t186 sky130_fd_pr__nfet_g5v0d10v5 ad=0.638 pd=4.69 as=0.638 ps=4.69 w=4.4 l=1
X322 DVSS.t137 D0.t1 sky130_fd_pr__diode_pw2nd_11v0 perim=3.16e+06 area=6.072e+11
X323 a_16261_n4916.t20 D93v3.t11 x3.R1.t75 VSS.t186 sky130_fd_pr__nfet_g5v0d10v5 ad=0.638 pd=4.69 as=0.638 ps=4.69 w=4.4 l=1
X324 x6.V1.t50 x9.V2.t37 VSS.t126 sky130_fd_pr__res_high_po_0p69 l=12.22
X325 x3.R1.t49 x8.V2.t49 VSS.t131 sky130_fd_pr__res_high_po_0p69 l=12.22
X326 x5.V2.t82 D43v3.t16 a_6164_n9984.t10 VSS.t243 sky130_fd_pr__nfet_g5v0d10v5 ad=0.638 pd=4.69 as=1.276 ps=9.38 w=4.4 l=1
X327 a_n1825_14638# a_n2121_15261# VDD.t192 VDD.t107 sky130_fd_pr__pfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.24375 ps=1.825 w=1.5 l=0.5
X328 DVSS.t110 a_n1825_4654# D33v3.t0 DVSS.t109 sky130_fd_pr__nfet_g5v0d10v5 ad=0.121875 pd=1.075 as=0.19875 ps=2.03 w=0.75 l=0.5
X329 DVDD.t39 a_n2559_n4073# a_n2603_n5122# DVDD.t38 sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.12 as=0.2478 ps=2.27 w=0.84 l=0.15
X330 ia_opamp_0.V2.t33 a_10431_n8604# VSS.t106 sky130_fd_pr__res_high_po_0p69 l=12.22
X331 VDD.t24 a_3421_764.t6 a_4215_764.t2 VDD.t23 sky130_fd_pr__pfet_g5v0d10v5 ad=4.35 pd=30.58 as=2.175 ps=15.29 w=15 l=1
X332 DVSS.t179 a_n2603_4862# a_n2577_4809# DVSS.t176 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.3975 ps=3.53 w=1.5 l=0.5
X333 a_n2577_n2679# a_n2603_n2626# DVSS.t142 DVSS.t138 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X334 x6.V1.t64 x9.V2.t46 VSS.t184 sky130_fd_pr__res_high_po_0p69 l=12.22
X335 x4.V2.t84 D43v3.t17 a_6164_n4916.t11 VSS.t243 sky130_fd_pr__nfet_g5v0d10v5 ad=0.638 pd=4.69 as=1.276 ps=9.38 w=4.4 l=1
X336 VOUT.t5 a_10431_n3536# VSS.t106 sky130_fd_pr__res_high_po_0p69 l=12.22
X337 x5.V2.t12 x4.V2.t13 VSS.t65 sky130_fd_pr__res_high_po_0p69 l=12.22
X338 DVSS.t174 a_n2603_14846# a_n2577_14793# DVSS.t170 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.3975 ps=3.53 w=1.5 l=0.5
X339 a_n2577_4809# a_n2603_4862# DVSS.t178 DVSS.t176 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X340 DVSS.t262 a_n2559_919# a_n2121_285# DVSS.t261 sky130_fd_pr__nfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.21 ps=1.78 w=1.5 l=0.5
X341 x6.V1.t86 x9.V2.t62 VSS.t64 sky130_fd_pr__res_high_po_0p69 l=12.22
X342 amp_biases_0.ibias3.t3 a_204_12823.t10 VDD.t38 VDD.t37 sky130_fd_pr__pfet_g5v0d10v5 ad=2.175 pd=15.29 as=2.175 ps=15.29 w=15 l=1
X343 VSS.t212 amp_biases_0.ibias4.t4 a_13231_764.t0 VSS.t211 sky130_fd_pr__nfet_g5v0d10v5 ad=4.4776 pd=31.46 as=4.4776 ps=31.46 w=15.44 l=1
X344 a_n1825_n7826# a_n2121_n7203# DVSS.t153 DVSS.t152 sky130_fd_pr__nfet_g5v0d10v5 ad=0.19875 pd=2.03 as=0.121875 ps=1.075 w=0.75 l=0.5
X345 x6.V1.t93 x9.V2.t69 VSS.t102 sky130_fd_pr__res_high_po_0p69 l=12.22
X346 AVOUT2.t16 a_3720_n9984.t11 VSS.t130 sky130_fd_pr__res_high_po_0p69 l=12.22
X347 DVSS.t185 a_n2603_n130# a_n2577_n183# DVSS.t182 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.3975 ps=3.53 w=1.5 l=0.5
X348 a_10431_n8604# VDD.t241 x6.V1.t53 VSS.t182 sky130_fd_pr__nfet_g5v0d10v5 ad=1.3833 pd=10.12 as=1.3833 ps=10.12 w=4.77 l=1
X349 a_3679_764.t1 x4.V2.t94 a_3421_764.t0 VSS.t90 sky130_fd_pr__nfet_g5v0d10v5 ad=4.785 pd=33.58 as=4.785 ps=33.58 w=16.5 l=1
X350 DVSS.t123 a_n2559_15895# a_n2121_15261# DVSS.t122 sky130_fd_pr__nfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.21 ps=1.78 w=1.5 l=0.5
X351 AVOUT1.t15 a_3720_n4916.t10 VSS.t130 sky130_fd_pr__res_high_po_0p69 l=12.22
X352 a_16951_764.t3 x6.V1.t94 a_16415_764.t2 VSS.t239 sky130_fd_pr__nfet_g5v0d10v5 ad=4.785 pd=33.58 as=4.785 ps=33.58 w=16.5 l=1
X353 a_n2559_n4073# D7.t1 DVSS.t51 DVSS.t50 sky130_fd_pr__nfet_01v8 ad=0.2478 pd=2.27 as=0.1176 ps=1.12 w=0.84 l=0.15
X354 a_10431_n3536# VDD.t242 x3.R1.t92 VSS.t182 sky130_fd_pr__nfet_g5v0d10v5 ad=1.3833 pd=10.12 as=1.3833 ps=10.12 w=4.77 l=1
X355 AVOUT1.t27 amp_biases_0.ibias1.t4 VSS.t205 VSS.t204 sky130_fd_pr__nfet_g5v0d10v5 ad=5.51 pd=38.58 as=5.51 ps=38.58 w=19 l=1
X356 x5.V2.t39 x4.V2.t39 VSS.t40 sky130_fd_pr__res_high_po_0p69 l=12.22
X357 a_16261_n9984.t22 D93v3.t12 x6.V1.t2 VSS.t11 sky130_fd_pr__nfet_g5v0d10v5 ad=1.276 pd=9.38 as=0.638 ps=4.69 w=4.4 l=1
X358 x6.V1.t30 x9.V2.t16 VSS.t131 sky130_fd_pr__res_high_po_0p69 l=12.22
X359 x3.R1.t17 x8.V2.t14 VSS.t79 sky130_fd_pr__res_high_po_0p69 l=12.22
X360 VDD.t40 a_204_12823.t11 amp_biases_0.ibias2.t3 VDD.t39 sky130_fd_pr__pfet_g5v0d10v5 ad=2.175 pd=15.29 as=2.175 ps=15.29 w=15 l=1
X361 x6.V1.t3 D93v3.t13 a_16261_n9984.t21 VSS.t12 sky130_fd_pr__nfet_g5v0d10v5 ad=0.638 pd=4.69 as=1.276 ps=9.38 w=4.4 l=1
X362 a_16261_n4916.t19 D93v3.t14 x3.R1.t74 VSS.t11 sky130_fd_pr__nfet_g5v0d10v5 ad=1.276 pd=9.38 as=0.638 ps=4.69 w=4.4 l=1
X363 a_n2577_n5175# a_n2603_n5122# DVSS.t130 DVSS.t126 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X364 AVOUT2.t21 a_3720_n9984.t12 VSS.t200 sky130_fd_pr__res_high_po_0p69 l=12.22
X365 a_n2577_7305# a_n2603_7358# DVSS.t232 DVSS.t229 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X366 VDD.t207 DVSS.t311 VDD.t206 VDD.t205 sky130_fd_pr__pfet_g5v0d10v5 ad=0.265 pd=2.53 as=0 ps=0 w=1 l=1
X367 x3.R1.t73 D93v3.t15 a_16261_n4916.t18 VSS.t12 sky130_fd_pr__nfet_g5v0d10v5 ad=0.638 pd=4.69 as=1.276 ps=9.38 w=4.4 l=1
X368 VOUT.t6 amp_biases_0.ibias5.t4 VSS.t110 VSS.t109 sky130_fd_pr__nfet_g5v0d10v5 ad=5.51 pd=38.58 as=5.51 ps=38.58 w=19 l=1
X369 ia_opamp_0.V2.t36 a_1031_764.t5 VDD.t231 VDD.t230 sky130_fd_pr__pfet_g5v0d10v5 ad=2.755 pd=19.29 as=5.51 ps=38.58 w=19 l=1
X370 DVSS.t56 D2.t1 sky130_fd_pr__diode_pw2nd_11v0 perim=3.16e+06 area=6.072e+11
X371 DVSS.t25 a_n2603_n10114# a_n2577_n10167# DVSS.t22 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.3975 ps=3.53 w=1.5 l=0.5
X372 VOUT.t32 a_16951_764.t5 VDD.t63 VDD.t62 sky130_fd_pr__pfet_g5v0d10v5 ad=2.755 pd=19.29 as=5.51 ps=38.58 w=19 l=1
X373 DVSS.t210 a_n2559_3415# a_n2121_2781# DVSS.t209 sky130_fd_pr__nfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.21 ps=1.78 w=1.5 l=0.5
X374 AVOUT1.t34 a_3720_n4916.t15 VSS.t200 sky130_fd_pr__res_high_po_0p69 l=12.22
X375 x5.V2.t22 x4.V2.t24 VSS.t51 sky130_fd_pr__res_high_po_0p69 l=12.22
X376 ia_opamp_0.V2.t30 a_13817_n9984.t15 VSS.t125 sky130_fd_pr__res_high_po_0p69 l=12.22
X377 a_3720_n9984.t5 D33v3.t12 x5.V2.t59 VSS.t195 sky130_fd_pr__nfet_g5v0d10v5 ad=0.6351 pd=4.67 as=0.6351 ps=4.67 w=4.38 l=1
X378 DVSS.t222 a_n2559_13399# a_n2121_12765# DVSS.t221 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.3975 ps=3.53 w=1.5 l=0.5
X379 VDD.t210 DVSS.t312 VDD.t209 VDD.t208 sky130_fd_pr__pfet_g5v0d10v5 ad=0.265 pd=2.53 as=0 ps=0 w=1 l=1
X380 VOUT.t11 a_13817_n4916.t2 VSS.t125 sky130_fd_pr__res_high_po_0p69 l=12.22
X381 x5.V2.t35 x4.V2.t33 VSS.t143 sky130_fd_pr__res_high_po_0p69 l=12.22
X382 a_n1825_12142# a_n2121_12765# DVSS.t107 DVSS.t106 sky130_fd_pr__nfet_g5v0d10v5 ad=0.19875 pd=2.03 as=0.121875 ps=1.075 w=0.75 l=0.5
X383 x3.R1.t29 x8.V2.t24 VSS.t65 sky130_fd_pr__res_high_po_0p69 l=12.22
X384 a_3720_n4916.t4 D33v3.t13 x4.V2.t62 VSS.t195 sky130_fd_pr__nfet_g5v0d10v5 ad=0.6351 pd=4.67 as=0.6351 ps=4.67 w=4.38 l=1
X385 DVSS.t283 VDD.t243 DVSS.t282 DVSS.t281 sky130_fd_pr__nfet_g5v0d10v5 ad=0.19875 pd=2.03 as=0 ps=0 w=0.75 l=1
X386 amp_biases_0.ibias2.t2 a_204_12823.t12 VDD.t75 VDD.t74 sky130_fd_pr__pfet_g5v0d10v5 ad=2.175 pd=15.29 as=2.175 ps=15.29 w=15 l=1
X387 DVSS.t280 VDD.t244 DVSS.t279 DVSS.t278 sky130_fd_pr__nfet_g5v0d10v5 ad=0.19875 pd=2.03 as=0 ps=0 w=0.75 l=1
X388 x3.R1.t50 x8.V2.t50 VSS.t180 sky130_fd_pr__res_high_po_0p69 l=12.22
X389 x6.V1.t21 x9.V2.t11 VSS.t79 sky130_fd_pr__res_high_po_0p69 l=12.22
X390 DVSS.t92 a_n2603_n7618# a_n2577_n7671# DVSS.t88 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.3975 ps=3.53 w=1.5 l=0.5
X391 x6.V1.t27 D93v3.t16 a_16261_n9984.t20 VSS.t111 sky130_fd_pr__nfet_g5v0d10v5 ad=0.638 pd=4.69 as=0.638 ps=4.69 w=4.4 l=1
X392 x5.V2.t72 x4.V2.t73 VSS.t174 sky130_fd_pr__res_high_po_0p69 l=12.22
X393 a_13817_n9984.t7 D83v3.t2 x6.V1.t60 VSS.t193 sky130_fd_pr__nfet_g5v0d10v5 ad=0.6351 pd=4.67 as=0.6351 ps=4.67 w=4.38 l=1
X394 x3.R1.t72 D93v3.t17 a_16261_n4916.t17 VSS.t111 sky130_fd_pr__nfet_g5v0d10v5 ad=0.638 pd=4.69 as=0.638 ps=4.69 w=4.4 l=1
X395 VDD.t174 a_237_764.t2 a_237_764.t3 VDD.t173 sky130_fd_pr__pfet_g5v0d10v5 ad=4.35 pd=30.58 as=2.175 ps=15.29 w=15 l=1
X396 DVSS.t132 D6.t0 sky130_fd_pr__diode_pw2nd_11v0 perim=3.16e+06 area=6.072e+11
X397 AVOUT2.t20 a_6164_n9984.t22 VSS.t183 sky130_fd_pr__res_high_po_0p69 l=12.22
X398 a_n1825_14638# a_n2121_15261# DVSS.t236 DVSS.t235 sky130_fd_pr__nfet_g5v0d10v5 ad=0.19875 pd=2.03 as=0.121875 ps=1.075 w=0.75 l=0.5
X399 a_n2121_2781# a_n2577_2313# VDD.t101 VDD.t100 sky130_fd_pr__pfet_g5v0d10v5 ad=0.2142 pd=1.99 as=0.2142 ps=1.99 w=0.42 l=1
X400 x6.V1.t84 x9.V2.t60 VSS.t65 sky130_fd_pr__res_high_po_0p69 l=12.22
X401 x3.R1.t89 x8.V2.t66 VSS.t145 sky130_fd_pr__res_high_po_0p69 l=12.22
X402 x6.V1.t5 D93v3.t18 a_16261_n9984.t19 VSS.t22 sky130_fd_pr__nfet_g5v0d10v5 ad=0.638 pd=4.69 as=0.638 ps=4.69 w=4.4 l=1
X403 a_13817_n4916.t12 D83v3.t3 x3.R1.t64 VSS.t193 sky130_fd_pr__nfet_g5v0d10v5 ad=0.6351 pd=4.67 as=0.6351 ps=4.67 w=4.38 l=1
X404 AVOUT1.t26 a_6164_n4916.t24 VSS.t183 sky130_fd_pr__res_high_po_0p69 l=12.22
X405 VSS.t83 amp_biases_0.ibias5.t5 a_16415_764.t0 VSS.t82 sky130_fd_pr__nfet_g5v0d10v5 ad=4.4776 pd=31.46 as=4.4776 ps=31.46 w=15.44 l=1
X406 VSS.t134 ia_opamp_0.ibias.t4 a_495_764.t1 VSS.t133 sky130_fd_pr__nfet_g5v0d10v5 ad=4.4776 pd=31.46 as=4.4776 ps=31.46 w=15.44 l=1
X407 DVSS.t31 a_n1825_7150# D23v3.t0 DVSS.t30 sky130_fd_pr__nfet_g5v0d10v5 ad=0.121875 pd=1.075 as=0.19875 ps=2.03 w=0.75 l=0.5
X408 x6.V1.t91 x9.V2.t67 VSS.t180 sky130_fd_pr__res_high_po_0p69 l=12.22
X409 x3.R1.t20 x8.V2.t16 VSS.t112 sky130_fd_pr__res_high_po_0p69 l=12.22
X410 x3.R1.t71 D93v3.t19 a_16261_n4916.t16 VSS.t22 sky130_fd_pr__nfet_g5v0d10v5 ad=0.638 pd=4.69 as=0.638 ps=4.69 w=4.4 l=1
X411 x5.V2.t36 D23v3.t4 a_2308_n9984.t2 VSS.t147 sky130_fd_pr__nfet_g5v0d10v5 ad=0.67425 pd=4.94 as=0.67425 ps=4.94 w=4.65 l=1
X412 ia_opamp_0.V2.t5 a_12405_n9984.t0 VSS.t58 sky130_fd_pr__res_high_po_0p69 l=12.22
X413 ia_opamp_0.V2.t1 a_16261_n9984.t1 VSS.t26 sky130_fd_pr__res_high_po_0p69 l=12.22
X414 x4.V2.t36 D23v3.t5 a_2308_n4916.t2 VSS.t147 sky130_fd_pr__nfet_g5v0d10v5 ad=0.67425 pd=4.94 as=0.67425 ps=4.94 w=4.65 l=1
X415 a_237_764.t1 a_237_764.t0 VDD.t172 VDD.t171 sky130_fd_pr__pfet_g5v0d10v5 ad=2.175 pd=15.29 as=4.35 ps=30.58 w=15 l=1
X416 x5.V2.t86 x4.V2.t87 VSS.t98 sky130_fd_pr__res_high_po_0p69 l=12.22
X417 VOUT.t16 a_12405_n4916.t2 VSS.t58 sky130_fd_pr__res_high_po_0p69 l=12.22
X418 a_n2559_n6569# D8.t0 DVSS.t20 DVSS.t19 sky130_fd_pr__nfet_01v8 ad=0.2478 pd=2.27 as=0.1176 ps=1.12 w=0.84 l=0.15
X419 x3.R1.t40 x8.V2.t39 VSS.t4 sky130_fd_pr__res_high_po_0p69 l=12.22
X420 VOUT.t22 a_16261_n4916.t10 VSS.t26 sky130_fd_pr__res_high_po_0p69 l=12.22
X421 a_n2121_2781# a_n2559_3415# DVSS.t208 DVSS.t207 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X422 DVSS.t206 a_n2559_3415# a_n2603_2366# DVSS.t205 sky130_fd_pr__nfet_01v8 ad=0.1176 pd=1.12 as=0.2478 ps=2.27 w=0.84 l=0.15
X423 VDD.t114 a_n1825_2158# D43v3.t1 VDD.t113 sky130_fd_pr__pfet_g5v0d10v5 ad=0.24375 pd=1.825 as=0.3975 ps=3.53 w=1.5 l=0.5
X424 x6.V1.t54 x9.V2.t40 VSS.t145 sky130_fd_pr__res_high_po_0p69 l=12.22
X425 x3.R1.t30 x8.V2.t25 VSS.t152 sky130_fd_pr__res_high_po_0p69 l=12.22
X426 x5.V2.t27 x4.V2.t26 VSS.t126 sky130_fd_pr__res_high_po_0p69 l=12.22
X427 a_n2577_n7671# a_n2603_n7618# DVSS.t91 DVSS.t88 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X428 x6.V1.t38 x9.V2.t25 VSS.t112 sky130_fd_pr__res_high_po_0p69 l=12.22
X429 x3.R1.t5 x8.V2.t5 VSS.t40 sky130_fd_pr__res_high_po_0p69 l=12.22
X430 x6.V1.t14 D73v3.t6 a_12405_n9984.t3 VSS.t52 sky130_fd_pr__nfet_g5v0d10v5 ad=0.67425 pd=4.94 as=0.67425 ps=4.94 w=4.65 l=1
X431 a_n2559_n9065# D9.t2 DVDD.t33 DVDD.t32 sky130_fd_pr__pfet_01v8_hvt ad=0.2478 pd=2.27 as=0.1176 ps=1.12 w=0.84 l=0.15
X432 x3.R1.t24 x8.V2.t20 VSS.t132 sky130_fd_pr__res_high_po_0p69 l=12.22
X433 a_16261_n9984.t18 D93v3.t20 x6.V1.t6 VSS.t1 sky130_fd_pr__nfet_g5v0d10v5 ad=0.638 pd=4.69 as=0.638 ps=4.69 w=4.4 l=1
X434 x3.R1.t8 D73v3.t7 a_12405_n4916.t4 VSS.t52 sky130_fd_pr__nfet_g5v0d10v5 ad=0.67425 pd=4.94 as=0.67425 ps=4.94 w=4.65 l=1
X435 a_16261_n4916.t15 D93v3.t21 x3.R1.t70 VSS.t1 sky130_fd_pr__nfet_g5v0d10v5 ad=0.638 pd=4.69 as=0.638 ps=4.69 w=4.4 l=1
X436 VDD.t148 a_10583_764.t6 x8.V2.t45 VDD.t147 sky130_fd_pr__pfet_g5v0d10v5 ad=2.755 pd=19.29 as=2.755 ps=19.29 w=19 l=1
X437 a_n2121_5277# a_n2559_5911# DVSS.t62 DVSS.t61 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X438 a_2308_n9984.t1 D23v3.t6 x5.V2.t23 VSS.t120 sky130_fd_pr__nfet_g5v0d10v5 ad=0.67425 pd=4.94 as=0.67425 ps=4.94 w=4.65 l=1
X439 DVSS.t60 a_n2559_5911# a_n2603_4862# DVSS.t59 sky130_fd_pr__nfet_01v8 ad=0.1176 pd=1.12 as=0.2478 ps=2.27 w=0.84 l=0.15
X440 VDD.t103 a_n1825_4654# D33v3.t1 VDD.t102 sky130_fd_pr__pfet_g5v0d10v5 ad=0.24375 pd=1.825 as=0.3975 ps=3.53 w=1.5 l=0.5
X441 x6.V1.t52 x9.V2.t39 VSS.t4 sky130_fd_pr__res_high_po_0p69 l=12.22
X442 AVOUT2.t31 a_6164_n9984.t26 VSS.t242 sky130_fd_pr__res_high_po_0p69 l=12.22
X443 a_16261_n9984.t17 D93v3.t22 x6.V1.t0 VSS.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=0.638 pd=4.69 as=0.638 ps=4.69 w=4.4 l=1
X444 a_3414_281.t1 a_4215_764.t1 sky130_fd_pr__cap_mim_m3_1 l=6.9 w=6.9
X445 AVOUT2.t32 a_6164_n9984.t27 VSS.t172 sky130_fd_pr__res_high_po_0p69 l=12.22
X446 a_2308_n4916.t1 D23v3.t7 x4.V2.t25 VSS.t120 sky130_fd_pr__nfet_g5v0d10v5 ad=0.67425 pd=4.94 as=0.67425 ps=4.94 w=4.65 l=1
X447 AVOUT1.t33 a_6164_n4916.t28 VSS.t242 sky130_fd_pr__res_high_po_0p69 l=12.22
X448 x5.V2.t53 x4.V2.t54 VSS.t100 sky130_fd_pr__res_high_po_0p69 l=12.22
X449 x6.V1.t56 x9.V2.t41 VSS.t152 sky130_fd_pr__res_high_po_0p69 l=12.22
X450 a_16261_n4916.t14 D93v3.t23 x3.R1.t69 VSS.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=0.638 pd=4.69 as=0.638 ps=4.69 w=4.4 l=1
X451 AVOUT1.t22 a_6164_n4916.t22 VSS.t172 sky130_fd_pr__res_high_po_0p69 l=12.22
X452 x9.V2.t45 amp_biases_0.ibias4.t5 VSS.t214 VSS.t213 sky130_fd_pr__nfet_g5v0d10v5 ad=5.51 pd=38.58 as=5.51 ps=38.58 w=19 l=1
X453 DVSS.t260 a_n2559_919# a_n2121_285# DVSS.t259 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X454 AVOUT2.t36 a_3720_n9984.t15 VSS.t153 sky130_fd_pr__res_high_po_0p69 l=12.22
X455 DVSS.t24 a_n2603_n10114# a_n2577_n10167# DVSS.t22 sky130_fd_pr__nfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.21 ps=1.78 w=1.5 l=0.5
X456 x6.V1.t90 x9.V2.t66 VSS.t40 sky130_fd_pr__res_high_po_0p69 l=12.22
X457 DVSS.t148 a_n2603_9854# a_n2577_9801# DVSS.t146 sky130_fd_pr__nfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.21 ps=1.78 w=1.5 l=0.5
X458 AVOUT1.t20 a_3720_n4916.t13 VSS.t153 sky130_fd_pr__res_high_po_0p69 l=12.22
X459 DVSS.t81 a_n2559_n1577# a_n2121_n2211# DVSS.t80 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X460 a_n2559_10903# D1.t2 DVDD.t9 DVDD.t8 sky130_fd_pr__pfet_01v8_hvt ad=0.2478 pd=2.27 as=0.1176 ps=1.12 w=0.84 l=0.15
X461 a_n2121_n7203# a_n2559_n6569# DVSS.t101 DVSS.t100 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X462 x6.V1.t81 x9.V2.t59 VSS.t132 sky130_fd_pr__res_high_po_0p69 l=12.22
X463 x5.V2.t90 x4.V2.t91 VSS.t62 sky130_fd_pr__res_high_po_0p69 l=12.22
X464 VSS.t207 amp_biases_0.ibias1.t5 a_3679_764.t0 VSS.t206 sky130_fd_pr__nfet_g5v0d10v5 ad=4.4776 pd=31.46 as=4.4776 ps=31.46 w=15.44 l=1
X465 a_13767_764.t3 AVOUT2.t38 a_13231_764.t2 VSS.t203 sky130_fd_pr__nfet_g5v0d10v5 ad=4.785 pd=33.58 as=4.785 ps=33.58 w=16.5 l=1
X466 ia_opamp_0.V2.t18 a_13817_n9984.t2 VSS.t128 sky130_fd_pr__res_high_po_0p69 l=12.22
X467 x3.R1.t3 x8.V2.t3 VSS.t24 sky130_fd_pr__res_high_po_0p69 l=12.22
X468 ia_opamp_0.V2.t13 a_16261_n9984.t8 VSS.t144 sky130_fd_pr__res_high_po_0p69 l=12.22
X469 ia_opamp_0.V2.t11 ia_opamp_0.ibias.t5 VSS.t136 VSS.t135 sky130_fd_pr__nfet_g5v0d10v5 ad=5.51 pd=38.58 as=5.51 ps=38.58 w=19 l=1
X470 VOUT.t12 a_13817_n4916.t3 VSS.t128 sky130_fd_pr__res_high_po_0p69 l=12.22
X471 DVSS.t240 a_n2603_2366# a_n2577_2313# DVSS.t237 sky130_fd_pr__nfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.21 ps=1.78 w=1.5 l=0.5
X472 x3.R1.t46 x8.V2.t44 VSS.t85 sky130_fd_pr__res_high_po_0p69 l=12.22
X473 VOUT.t34 a_16261_n4916.t28 VSS.t144 sky130_fd_pr__res_high_po_0p69 l=12.22
X474 DVSS.t199 a_n2603_12350# a_n2577_12297# DVSS.t196 sky130_fd_pr__nfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.21 ps=1.78 w=1.5 l=0.5
X475 DVDD.t41 a_n2559_919# a_n2603_n130# DVDD.t40 sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.12 as=0.2478 ps=2.27 w=0.84 l=0.15
X476 x3.R1.t37 x8.V2.t36 VSS.t35 sky130_fd_pr__res_high_po_0p69 l=12.22
X477 AVOUT2.t7 a_2308_n9984.t4 VSS.t71 sky130_fd_pr__res_high_po_0p69 l=12.22
X478 AVOUT1.t10 a_2308_n4916.t4 VSS.t71 sky130_fd_pr__res_high_po_0p69 l=12.22
X479 a_n1825_n10322# a_n2121_n9699# DVSS.t6 DVSS.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=0.19875 pd=2.03 as=0.121875 ps=1.075 w=0.75 l=0.5
X480 x6.V1.t87 x9.V2.t63 VSS.t24 sky130_fd_pr__res_high_po_0p69 l=12.22
X481 x6.V1.t19 x9.V2.t9 VSS.t85 sky130_fd_pr__res_high_po_0p69 l=12.22
X482 x5.V2.t68 x4.V2.t69 VSS.t160 sky130_fd_pr__res_high_po_0p69 l=12.22
X483 VSS.t166 amp_biases_0.ibias3.t4 a_10047_764.t1 VSS.t165 sky130_fd_pr__nfet_g5v0d10v5 ad=4.4776 pd=31.46 as=4.4776 ps=31.46 w=15.44 l=1
X484 ia_opamp_0.V2.t31 a_12405_n9984.t7 VSS.t209 sky130_fd_pr__res_high_po_0p69 l=12.22
X485 x5.V2.t88 x4.V2.t89 VSS.t158 sky130_fd_pr__res_high_po_0p69 l=12.22
X486 VDD.t176 a_13767_764.t4 x9.V2.t54 VDD.t175 sky130_fd_pr__pfet_g5v0d10v5 ad=2.755 pd=19.29 as=2.755 ps=19.29 w=19 l=1
X487 VOUT.t26 a_12405_n4916.t7 VSS.t209 sky130_fd_pr__res_high_po_0p69 l=12.22
X488 x6.V1.t9 x9.V2.t3 VSS.t35 sky130_fd_pr__res_high_po_0p69 l=12.22
X489 VDD.t42 a_n1825_7150# D23v3.t1 VDD.t41 sky130_fd_pr__pfet_g5v0d10v5 ad=0.24375 pd=1.825 as=0.3975 ps=3.53 w=1.5 l=0.5
X490 x3.R1.t91 x8.V2.t68 VSS.t104 sky130_fd_pr__res_high_po_0p69 l=12.22
X491 ia_opamp_0.V2.t9 a_12405_n9984.t1 VSS.t101 sky130_fd_pr__res_high_po_0p69 l=12.22
X492 DVSS.t14 a_n2559_10903# a_n2121_10269# DVSS.t13 sky130_fd_pr__nfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.21 ps=1.78 w=1.5 l=0.5
X493 x3.R1.t93 x8.V2.t69 VSS.t42 sky130_fd_pr__res_high_po_0p69 l=12.22
X494 VOUT.t8 a_12405_n4916.t1 VSS.t101 sky130_fd_pr__res_high_po_0p69 l=12.22
X495 x5.V2.t85 x4.V2.t86 VSS.t30 sky130_fd_pr__res_high_po_0p69 l=12.22
X496 a_13817_n9984.t13 D83v3.t4 x6.V1.t77 VSS.t234 sky130_fd_pr__nfet_g5v0d10v5 ad=0.6351 pd=4.67 as=0.6351 ps=4.67 w=4.38 l=1
X497 VDD.t189 a_n1825_n5330# D73v3.t1 VDD.t188 sky130_fd_pr__pfet_g5v0d10v5 ad=0.24375 pd=1.825 as=0.3975 ps=3.53 w=1.5 l=0.5
X498 x5.V2.t2 x4.V2.t2 VSS.t5 sky130_fd_pr__res_high_po_0p69 l=12.22
X499 a_n2121_10269# a_n2559_10903# DVSS.t12 DVSS.t11 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X500 x3.R1.t88 x8.V2.t65 VSS.t157 sky130_fd_pr__res_high_po_0p69 l=12.22
X501 a_13817_n4916.t13 D83v3.t5 x3.R1.t65 VSS.t234 sky130_fd_pr__nfet_g5v0d10v5 ad=0.6351 pd=4.67 as=0.6351 ps=4.67 w=4.38 l=1
X502 x9.V2.t55 a_13767_764.t5 VDD.t178 VDD.t177 sky130_fd_pr__pfet_g5v0d10v5 ad=2.755 pd=19.29 as=5.51 ps=38.58 w=19 l=1
X503 x5.V2.t19 x4.V2.t20 VSS.t102 sky130_fd_pr__res_high_po_0p69 l=12.22
X504 a_n2577_n5175# a_n2121_n4707# VDD.t224 VDD.t223 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1365 pd=1.49 as=0.1113 ps=1.37 w=0.42 l=1
X505 a_n2577_2313# a_n2603_2366# DVSS.t239 DVSS.t237 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X506 a_n2559_13399# D0.t2 DVDD.t29 DVDD.t28 sky130_fd_pr__pfet_01v8_hvt ad=0.2478 pd=2.27 as=0.1176 ps=1.12 w=0.84 l=0.15
X507 DVSS.t32 D4.t1 sky130_fd_pr__diode_pw2nd_11v0 perim=3.16e+06 area=6.072e+11
X508 a_n2121_n9699# a_n2559_n9065# DVSS.t163 DVSS.t162 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X509 a_n2577_12297# a_n2603_12350# DVSS.t198 DVSS.t196 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X510 x6.V1.t26 x9.V2.t14 VSS.t104 sky130_fd_pr__res_high_po_0p69 l=12.22
X511 x5.V2.t76 x4.V2.t78 VSS.t59 sky130_fd_pr__res_high_po_0p69 l=12.22
X512 x6.V1.t10 x9.V2.t4 VSS.t42 sky130_fd_pr__res_high_po_0p69 l=12.22
X513 x5.V2.t37 x4.V2.t37 VSS.t150 sky130_fd_pr__res_high_po_0p69 l=12.22
X514 a_n2121_12765# a_n2559_13399# DVSS.t220 DVSS.t219 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X515 DVSS.t277 VDD.t245 DVSS.t276 DVSS.t275 sky130_fd_pr__nfet_g5v0d10v5 ad=0.19875 pd=2.03 as=0 ps=0 w=0.75 l=1
X516 VDD.t85 a_n1825_n7826# D83v3.t1 VDD.t84 sky130_fd_pr__pfet_g5v0d10v5 ad=0.24375 pd=1.825 as=0.3975 ps=3.53 w=1.5 l=0.5
X517 a_6164_n9984.t9 D43v3.t18 x5.V2.t77 VSS.t232 sky130_fd_pr__nfet_g5v0d10v5 ad=1.276 pd=9.38 as=0.638 ps=4.69 w=4.4 l=1
X518 DVSS.t173 a_n2603_14846# a_n2577_14793# DVSS.t170 sky130_fd_pr__nfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.21 ps=1.78 w=1.5 l=0.5
X519 x6.V1.t39 x9.V2.t26 VSS.t157 sky130_fd_pr__res_high_po_0p69 l=12.22
X520 a_16415_764.t1 x3.R1.t94 a_16157_764.t4 VSS.t96 sky130_fd_pr__nfet_g5v0d10v5 ad=4.785 pd=33.58 as=4.785 ps=33.58 w=16.5 l=1
X521 a_2564_12836# sky130_fd_sc_hvl__lsbuflv2hv_1_0[10].X.t3 a_204_12823.t0 VSS.t169 sky130_fd_pr__nfet_g5v0d10v5 ad=2.2388 pd=15.73 as=4.4776 ps=31.46 w=15.44 l=1
X522 a_n2577_n2679# a_n2121_n2211# VDD.t87 VDD.t86 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1365 pd=1.49 as=0.1113 ps=1.37 w=0.42 l=1
X523 a_6164_n4916.t10 D43v3.t19 x4.V2.t79 VSS.t232 sky130_fd_pr__nfet_g5v0d10v5 ad=1.276 pd=9.38 as=0.638 ps=4.69 w=4.4 l=1
X524 VDD.t213 DVSS.t313 VDD.t212 VDD.t211 sky130_fd_pr__pfet_g5v0d10v5 ad=0.265 pd=2.53 as=0 ps=0 w=1 l=1
X525 a_n2559_15895# ena.t2 DVDD.t43 DVDD.t42 sky130_fd_pr__pfet_01v8_hvt ad=0.2478 pd=2.27 as=0.1176 ps=1.12 w=0.84 l=0.15
X526 DVSS.t71 D3.t1 sky130_fd_pr__diode_pw2nd_11v0 perim=3.16e+06 area=6.072e+11
X527 DVSS.t141 a_n2603_n2626# a_n2577_n2679# DVSS.t138 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.3975 ps=3.53 w=1.5 l=0.5
X528 x9.V2.t49 a_13767_764.t6 VDD.t168 VDD.t167 sky130_fd_pr__pfet_g5v0d10v5 ad=2.755 pd=19.29 as=2.755 ps=19.29 w=19 l=1
X529 x5.V2.t49 x4.V2.t50 VSS.t180 sky130_fd_pr__res_high_po_0p69 l=12.22
X530 a_10583_764.t3 AVOUT1.t38 a_10047_764.t2 VSS.t78 sky130_fd_pr__nfet_g5v0d10v5 ad=4.785 pd=33.58 as=4.785 ps=33.58 w=16.5 l=1
X531 AVOUT2.t24 a_7399_764.t5 VDD.t146 VDD.t145 sky130_fd_pr__pfet_g5v0d10v5 ad=2.755 pd=19.29 as=5.51 ps=38.58 w=19 l=1
X532 a_n2121_15261# a_n2559_15895# DVSS.t121 DVSS.t120 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X533 x3.R1.t32 x8.V2.t27 VSS.t77 sky130_fd_pr__res_high_po_0p69 l=12.22
X534 ia_opamp_0.V2.t6 a_16261_n9984.t5 VSS.t66 sky130_fd_pr__res_high_po_0p69 l=12.22
X535 a_2308_n9984.t0 D23v3.t8 x5.V2.t24 VSS.t121 sky130_fd_pr__nfet_g5v0d10v5 ad=1.3485 pd=9.88 as=0.67425 ps=4.94 w=4.65 l=1
X536 VOUT.t18 a_16261_n4916.t6 VSS.t66 sky130_fd_pr__res_high_po_0p69 l=12.22
X537 DVSS.t10 a_n2559_10903# a_n2603_9854# DVSS.t9 sky130_fd_pr__nfet_01v8 ad=0.1176 pd=1.12 as=0.2478 ps=2.27 w=0.84 l=0.15
X538 a_2308_n4916.t0 D23v3.t9 x4.V2.t34 VSS.t121 sky130_fd_pr__nfet_g5v0d10v5 ad=1.3485 pd=9.88 as=0.67425 ps=4.94 w=4.65 l=1
X539 DVSS.t197 a_n2603_12350# a_n2577_12297# DVSS.t196 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.3975 ps=3.53 w=1.5 l=0.5
X540 x8.V2.t30 amp_biases_0.ibias3.t5 VSS.t168 VSS.t167 sky130_fd_pr__nfet_g5v0d10v5 ad=5.51 pd=38.58 as=5.51 ps=38.58 w=19 l=1
X541 x3.R1.t0 x8.V2.t0 VSS.t5 sky130_fd_pr__res_high_po_0p69 l=12.22
X542 a_n2577_2313# a_n2121_2781# VDD.t180 VDD.t179 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1365 pd=1.49 as=0.1113 ps=1.37 w=0.42 l=1
X543 x6.V1.t22 D93v3.t24 a_16261_n9984.t16 VSS.t97 sky130_fd_pr__nfet_g5v0d10v5 ad=0.638 pd=4.69 as=0.638 ps=4.69 w=4.4 l=1
X544 a_n2559_n1577# D6.t1 DVSS.t134 DVSS.t133 sky130_fd_pr__nfet_01v8 ad=0.2478 pd=2.27 as=0.1176 ps=1.12 w=0.84 l=0.15
X545 x3.R1.t85 x8.V2.t62 VSS.t38 sky130_fd_pr__res_high_po_0p69 l=12.22
X546 x5.V2.t78 D43v3.t20 a_6164_n9984.t8 VSS.t222 sky130_fd_pr__nfet_g5v0d10v5 ad=0.638 pd=4.69 as=0.638 ps=4.69 w=4.4 l=1
X547 x3.R1.t68 D93v3.t25 a_16261_n4916.t25 VSS.t97 sky130_fd_pr__nfet_g5v0d10v5 ad=0.638 pd=4.69 as=0.638 ps=4.69 w=4.4 l=1
X548 DVSS.t228 a_n1825_n5330# D73v3.t0 DVSS.t227 sky130_fd_pr__nfet_g5v0d10v5 ad=0.121875 pd=1.075 as=0.19875 ps=2.03 w=0.75 l=0.5
X549 DVSS.t218 a_n2559_13399# a_n2603_12350# DVSS.t217 sky130_fd_pr__nfet_01v8 ad=0.1176 pd=1.12 as=0.2478 ps=2.27 w=0.84 l=0.15
X550 AVOUT2.t13 a_6164_n9984.t19 VSS.t72 sky130_fd_pr__res_high_po_0p69 l=12.22
X551 x4.V2.t76 D43v3.t21 a_6164_n4916.t9 VSS.t222 sky130_fd_pr__nfet_g5v0d10v5 ad=0.638 pd=4.69 as=0.638 ps=4.69 w=4.4 l=1
X552 x6.V1.t72 x9.V2.t53 VSS.t77 sky130_fd_pr__res_high_po_0p69 l=12.22
X553 amp_biases_0.ibias4.t3 a_204_12823.t13 VDD.t77 VDD.t76 sky130_fd_pr__pfet_g5v0d10v5 ad=2.175 pd=15.29 as=2.175 ps=15.29 w=15 l=1
X554 AVOUT2.t15 a_334_n8604# VSS.t163 sky130_fd_pr__res_high_po_0p69 l=12.22
X555 AVOUT1.t8 a_6164_n4916.t4 VSS.t72 sky130_fd_pr__res_high_po_0p69 l=12.22
X556 a_n2577_n7671# a_n2121_n7203# VDD.t124 VDD.t123 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1365 pd=1.49 as=0.1113 ps=1.37 w=0.42 l=1
X557 x5.V2.t75 D43v3.t22 a_6164_n9984.t7 VSS.t223 sky130_fd_pr__nfet_g5v0d10v5 ad=0.638 pd=4.69 as=0.638 ps=4.69 w=4.4 l=1
X558 a_12405_n9984.t2 D73v3.t8 x6.V1.t15 VSS.t53 sky130_fd_pr__nfet_g5v0d10v5 ad=1.3485 pd=9.88 as=0.67425 ps=4.94 w=4.65 l=1
X559 a_12405_n4916.t3 D73v3.t9 x3.R1.t18 VSS.t53 sky130_fd_pr__nfet_g5v0d10v5 ad=1.3485 pd=9.88 as=0.67425 ps=4.94 w=4.65 l=1
X560 x4.V2.t77 D43v3.t23 a_6164_n4916.t8 VSS.t223 sky130_fd_pr__nfet_g5v0d10v5 ad=0.638 pd=4.69 as=0.638 ps=4.69 w=4.4 l=1
X561 AVOUT1.t23 a_334_n3536# VSS.t163 sky130_fd_pr__res_high_po_0p69 l=12.22
X562 a_n2577_14793# a_n2603_14846# DVSS.t172 DVSS.t170 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X563 a_n1825_4654# a_n2121_5277# DVSS.t244 DVSS.t243 sky130_fd_pr__nfet_g5v0d10v5 ad=0.19875 pd=2.03 as=0.121875 ps=1.075 w=0.75 l=0.5
X564 DVSS.t258 a_n2559_919# a_n2603_n130# DVSS.t257 sky130_fd_pr__nfet_01v8 ad=0.1176 pd=1.12 as=0.2478 ps=2.27 w=0.84 l=0.15
X565 a_n2559_n4073# D7.t2 DVDD.t15 DVDD.t14 sky130_fd_pr__pfet_01v8_hvt ad=0.2478 pd=2.27 as=0.1176 ps=1.12 w=0.84 l=0.15
X566 x6.V1.t51 x9.V2.t38 VSS.t5 sky130_fd_pr__res_high_po_0p69 l=12.22
X567 a_334_n8604# VDD.t246 x5.V2.t92 VSS.t23 sky130_fd_pr__nfet_g5v0d10v5 ad=1.3833 pd=10.12 as=1.3833 ps=10.12 w=4.77 l=1
X568 AVOUT2.t14 a_2308_n9984.t5 VSS.t162 sky130_fd_pr__res_high_po_0p69 l=12.22
X569 x5.V2.t40 D13v3.t4 a_1412_n9984# VSS.t155 sky130_fd_pr__nfet_g5v0d10v5 ad=0.70615 pd=5.16 as=1.4123 ps=10.32 w=4.87 l=1
X570 AVOUT2.t26 a_6164_n9984.t24 VSS.t28 sky130_fd_pr__res_high_po_0p69 l=12.22
X571 AVOUT1.t36 a_2308_n4916.t7 VSS.t162 sky130_fd_pr__res_high_po_0p69 l=12.22
X572 x6.V1.t92 x9.V2.t68 VSS.t38 sky130_fd_pr__res_high_po_0p69 l=12.22
X573 x4.V2.t41 D13v3.t5 a_1412_n4916# VSS.t155 sky130_fd_pr__nfet_g5v0d10v5 ad=0.70615 pd=5.16 as=1.4123 ps=10.32 w=4.87 l=1
X574 a_334_n3536# VDD.t247 x4.V2.t92 VSS.t23 sky130_fd_pr__nfet_g5v0d10v5 ad=1.3833 pd=10.12 as=1.3833 ps=10.12 w=4.77 l=1
X575 AVOUT1.t1 a_6164_n4916.t1 VSS.t28 sky130_fd_pr__res_high_po_0p69 l=12.22
X576 VDD.t79 a_204_12823.t14 amp_biases_0.ibias3.t2 VDD.t78 sky130_fd_pr__pfet_g5v0d10v5 ad=2.175 pd=15.29 as=2.175 ps=15.29 w=15 l=1
X577 DVSS.t58 a_n2559_5911# a_n2121_5277# DVSS.t57 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X578 DVSS.t73 a_n1825_n7826# D83v3.t0 DVSS.t72 sky130_fd_pr__nfet_g5v0d10v5 ad=0.121875 pd=1.075 as=0.19875 ps=2.03 w=0.75 l=0.5
X579 x5.V2.t28 x4.V2.t27 VSS.t104 sky130_fd_pr__res_high_po_0p69 l=12.22
X580 DVSS.t117 a_n2559_15895# a_n2603_14846# DVSS.t116 sky130_fd_pr__nfet_01v8 ad=0.1176 pd=1.12 as=0.2478 ps=2.27 w=0.84 l=0.15
X581 ia_opamp_0.V2.t29 a_16261_n9984.t28 VSS.t181 sky130_fd_pr__res_high_po_0p69 l=12.22
X582 x5.V2.t89 x4.V2.t90 VSS.t217 sky130_fd_pr__res_high_po_0p69 l=12.22
X583 VOUT.t21 a_16261_n4916.t9 VSS.t181 sky130_fd_pr__res_high_po_0p69 l=12.22
X584 a_n2577_n10167# a_n2121_n9699# VDD.t13 VDD.t12 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1365 pd=1.49 as=0.1113 ps=1.37 w=0.42 l=1
X585 a_9782_281.t0 x8.V2.t32 VSS.t173 sky130_fd_pr__res_high_po_0p69 l=3.2
X586 DVSS.t129 a_n2603_n5122# a_n2577_n5175# DVSS.t126 sky130_fd_pr__nfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.21 ps=1.78 w=1.5 l=0.5
X587 DVSS.t184 a_n2603_n130# a_n2577_n183# DVSS.t182 sky130_fd_pr__nfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.21 ps=1.78 w=1.5 l=0.5
X588 DVSS.t128 a_n2603_n5122# a_n2577_n5175# DVSS.t126 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.3975 ps=3.53 w=1.5 l=0.5
X589 x5.V2.t60 D33v3.t14 a_3720_n9984.t4 VSS.t88 sky130_fd_pr__nfet_g5v0d10v5 ad=0.6351 pd=4.67 as=0.6351 ps=4.67 w=4.38 l=1
X590 x3.R1.t36 x8.V2.t33 VSS.t164 sky130_fd_pr__res_high_po_0p69 l=12.22
X591 x5.V2.t15 x4.V2.t16 VSS.t77 sky130_fd_pr__res_high_po_0p69 l=12.22
X592 a_6164_n9984.t6 D43v3.t24 x5.V2.t9 VSS.t54 sky130_fd_pr__nfet_g5v0d10v5 ad=0.638 pd=4.69 as=0.638 ps=4.69 w=4.4 l=1
X593 a_n2121_n2211# a_n2559_n1577# DVSS.t79 DVSS.t78 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X594 x3.R1.t45 x8.V2.t43 VSS.t27 sky130_fd_pr__res_high_po_0p69 l=12.22
X595 x6.V1.t69 D63v3.t4 a_11509_n9984# VSS.t221 sky130_fd_pr__nfet_g5v0d10v5 ad=0.70615 pd=5.16 as=1.4123 ps=10.32 w=4.87 l=1
X596 x4.V2.t18 D33v3.t15 a_3720_n4916.t3 VSS.t88 sky130_fd_pr__nfet_g5v0d10v5 ad=0.6351 pd=4.67 as=0.6351 ps=4.67 w=4.38 l=1
X597 x5.V2.t54 x4.V2.t55 VSS.t177 sky130_fd_pr__res_high_po_0p69 l=12.22
X598 x3.R1.t10 x8.V2.t9 VSS.t59 sky130_fd_pr__res_high_po_0p69 l=12.22
X599 x3.R1.t56 D63v3.t5 a_11509_n4916# VSS.t221 sky130_fd_pr__nfet_g5v0d10v5 ad=0.70615 pd=5.16 as=1.4123 ps=10.32 w=4.87 l=1
X600 a_6164_n4916.t7 D43v3.t25 x4.V2.t11 VSS.t54 sky130_fd_pr__nfet_g5v0d10v5 ad=0.638 pd=4.69 as=0.638 ps=4.69 w=4.4 l=1
X601 a_13231_764.t1 x9.V2.t70 a_12973_764.t4 VSS.t240 sky130_fd_pr__nfet_g5v0d10v5 ad=4.785 pd=33.58 as=4.785 ps=33.58 w=16.5 l=1
X602 a_n2121_7773# a_n2559_8407# DVSS.t39 DVSS.t38 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X603 VDD.t229 a_1031_764.t6 ia_opamp_0.V2.t35 VDD.t228 sky130_fd_pr__pfet_g5v0d10v5 ad=2.755 pd=19.29 as=2.755 ps=19.29 w=19 l=1
X604 amp_biases_0.ibias5.t1 amp_biases_0.ibias5.t0 VSS.t189 VSS.t188 sky130_fd_pr__nfet_g5v0d10v5 ad=4.4776 pd=31.46 as=4.4776 ps=31.46 w=15.44 l=1
X605 VDD.t65 a_16951_764.t6 VOUT.t31 VDD.t64 sky130_fd_pr__pfet_g5v0d10v5 ad=2.755 pd=19.29 as=2.755 ps=19.29 w=19 l=1
X606 a_n2577_n183# a_n2121_285# VDD.t56 VDD.t55 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1365 pd=1.49 as=0.1113 ps=1.37 w=0.42 l=1
X607 AVOUT2.t22 a_3720_n9984.t13 VSS.t151 sky130_fd_pr__res_high_po_0p69 l=12.22
X608 a_n2577_4809# a_n2121_5277# VDD.t197 VDD.t196 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1365 pd=1.49 as=0.1113 ps=1.37 w=0.42 l=1
X609 DVSS.t90 a_n2603_n7618# a_n2577_n7671# DVSS.t88 sky130_fd_pr__nfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.21 ps=1.78 w=1.5 l=0.5
X610 x5.V2.t52 x4.V2.t53 VSS.t184 sky130_fd_pr__res_high_po_0p69 l=12.22
X611 DVSS.t140 a_n2603_n2626# a_n2577_n2679# DVSS.t138 sky130_fd_pr__nfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.21 ps=1.78 w=1.5 l=0.5
X612 x5.V2.t50 x4.V2.t51 VSS.t131 sky130_fd_pr__res_high_po_0p69 l=12.22
X613 a_n2577_n7671# a_n2603_n7618# DVSS.t89 DVSS.t88 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X614 AVOUT1.t19 a_3720_n4916.t12 VSS.t151 sky130_fd_pr__res_high_po_0p69 l=12.22
X615 x5.V2.t67 x4.V2.t68 VSS.t27 sky130_fd_pr__res_high_po_0p69 l=12.22
X616 x6.V1.t58 D83v3.t6 a_13817_n9984.t5 VSS.t190 sky130_fd_pr__nfet_g5v0d10v5 ad=0.6351 pd=4.67 as=0.6351 ps=4.67 w=4.38 l=1
X617 x6.V1.t45 x9.V2.t32 VSS.t164 sky130_fd_pr__res_high_po_0p69 l=12.22
X618 x6.V1.t7 x9.V2.t1 VSS.t27 sky130_fd_pr__res_high_po_0p69 l=12.22
X619 DVSS.t250 a_n2559_n4073# a_n2121_n4707# DVSS.t249 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.3975 ps=3.53 w=1.5 l=0.5
X620 a_10959_n8604# D53v3.t2 x6.V1.t29 VSS.t119 sky130_fd_pr__nfet_g5v0d10v5 ad=1.3833 pd=10.12 as=1.3833 ps=10.12 w=4.77 l=1
X621 x3.R1.t42 D83v3.t7 a_13817_n4916.t5 VSS.t190 sky130_fd_pr__nfet_g5v0d10v5 ad=0.6351 pd=4.67 as=0.6351 ps=4.67 w=4.38 l=1
X622 x6.V1.t47 x9.V2.t34 VSS.t59 sky130_fd_pr__res_high_po_0p69 l=12.22
X623 x3.R1.t27 x8.V2.t22 VSS.t60 sky130_fd_pr__res_high_po_0p69 l=12.22
X624 ia_opamp_0.V2.t0 a_16261_n9984.t0 VSS.t25 sky130_fd_pr__res_high_po_0p69 l=12.22
X625 a_16261_n9984.t15 D93v3.t26 x6.V1.t23 VSS.t20 sky130_fd_pr__nfet_g5v0d10v5 ad=0.638 pd=4.69 as=0.638 ps=4.69 w=4.4 l=1
X626 VDD.t116 a_204_12823.t1 a_204_12823.t2 VDD.t115 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=1
X627 x6.V1.t59 D83v3.t8 a_13817_n9984.t6 VSS.t191 sky130_fd_pr__nfet_g5v0d10v5 ad=0.6351 pd=4.67 as=1.2702 ps=9.34 w=4.38 l=1
X628 AVOUT2.t8 a_3720_n9984.t2 VSS.t80 sky130_fd_pr__res_high_po_0p69 l=12.22
X629 a_16261_n4916.t24 D93v3.t27 x3.R1.t67 VSS.t20 sky130_fd_pr__nfet_g5v0d10v5 ad=0.638 pd=4.69 as=0.638 ps=4.69 w=4.4 l=1
X630 a_10959_n3536# D53v3.t3 x3.R1.t26 VSS.t119 sky130_fd_pr__nfet_g5v0d10v5 ad=1.3833 pd=10.12 as=1.3833 ps=10.12 w=4.77 l=1
X631 VOUT.t19 a_16261_n4916.t7 VSS.t25 sky130_fd_pr__res_high_po_0p69 l=12.22
X632 VDD.t71 a_4215_764.t4 AVOUT1.t12 VDD.t70 sky130_fd_pr__pfet_g5v0d10v5 ad=5.51 pd=38.58 as=2.755 ps=19.29 w=19 l=1
X633 x3.R1.t62 D83v3.t9 a_13817_n4916.t10 VSS.t191 sky130_fd_pr__nfet_g5v0d10v5 ad=0.6351 pd=4.67 as=1.2702 ps=9.34 w=4.38 l=1
X634 a_n1825_7150# a_n2121_7773# DVSS.t189 DVSS.t188 sky130_fd_pr__nfet_g5v0d10v5 ad=0.19875 pd=2.03 as=0.121875 ps=1.075 w=0.75 l=0.5
X635 AVOUT1.t16 a_3720_n4916.t11 VSS.t80 sky130_fd_pr__res_high_po_0p69 l=12.22
X636 a_n2577_7305# a_n2121_7773# VDD.t153 VDD.t152 sky130_fd_pr__pfet_g5v0d10v5 ad=0.1365 pd=1.49 as=0.1113 ps=1.37 w=0.42 l=1
X637 a_n2559_n6569# D8.t1 DVDD.t3 DVDD.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.2478 pd=2.27 as=0.1176 ps=1.12 w=0.84 l=0.15
X638 ia_opamp_0.V2.t27 a_13817_n9984.t14 VSS.t245 sky130_fd_pr__res_high_po_0p69 l=12.22
X639 x5.V2.t45 x4.V2.t47 VSS.t6 sky130_fd_pr__res_high_po_0p69 l=12.22
X640 a_n2577_n10167# a_n2603_n10114# DVSS.t23 DVSS.t22 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X641 VDD.t108 a_n1825_14638# sky130_fd_sc_hvl__lsbuflv2hv_1_0[10].X.t1 VDD.t107 sky130_fd_pr__pfet_g5v0d10v5 ad=0.24375 pd=1.825 as=0.3975 ps=3.53 w=1.5 l=0.5
X642 x3.R1.t21 x8.V2.t17 VSS.t114 sky130_fd_pr__res_high_po_0p69 l=12.22
X643 ia_opamp_0.V2.t32 a_16261_n9984.t29 VSS.t246 sky130_fd_pr__res_high_po_0p69 l=12.22
X644 VOUT.t35 a_13817_n4916.t14 VSS.t245 sky130_fd_pr__res_high_po_0p69 l=12.22
X645 DVSS.t37 a_n2559_8407# a_n2121_7773# DVSS.t36 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X646 VOUT.t36 a_16261_n4916.t29 VSS.t246 sky130_fd_pr__res_high_po_0p69 l=12.22
X647 AVOUT1.t13 a_4215_764.t5 VDD.t73 VDD.t72 sky130_fd_pr__pfet_g5v0d10v5 ad=2.755 pd=19.29 as=2.755 ps=19.29 w=19 l=1
X648 DVSS.t99 a_n2559_n6569# a_n2121_n7203# DVSS.t98 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.3975 ps=3.53 w=1.5 l=0.5
X649 DVSS.t77 a_n2559_n1577# a_n2121_n2211# DVSS.t76 sky130_fd_pr__nfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.21 ps=1.78 w=1.5 l=0.5
X650 x6.V1.t89 x9.V2.t65 VSS.t60 sky130_fd_pr__res_high_po_0p69 l=12.22
X651 AVOUT2.t6 amp_biases_0.ibias2.t5 VSS.t70 VSS.t69 sky130_fd_pr__nfet_g5v0d10v5 ad=5.51 pd=38.58 as=5.51 ps=38.58 w=19 l=1
X652 DVSS.t8 a_n2559_10903# a_n2121_10269# DVSS.t7 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X653 a_n1825_9646# a_n2121_10269# DVSS.t155 DVSS.t154 sky130_fd_pr__nfet_g5v0d10v5 ad=0.19875 pd=2.03 as=0.121875 ps=1.075 w=0.75 l=0.5
X654 AVOUT2.t37 a_2308_n9984.t7 VSS.t127 sky130_fd_pr__res_high_po_0p69 l=12.22
X655 DVSS.t238 a_n2603_2366# a_n2577_2313# DVSS.t237 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X656 a_n2121_n4707# a_n2559_n4073# DVSS.t248 DVSS.t247 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X657 a_862_n8604# D03v3.t2 x5.V2.t34 VSS.t146 sky130_fd_pr__nfet_g5v0d10v5 ad=1.3833 pd=10.12 as=1.3833 ps=10.12 w=4.77 l=1
X658 AVOUT2.t35 a_6164_n9984.t29 VSS.t210 sky130_fd_pr__res_high_po_0p69 l=12.22
X659 VDD.t20 a_4215_764.t6 AVOUT1.t6 VDD.t19 sky130_fd_pr__pfet_g5v0d10v5 ad=2.755 pd=19.29 as=2.755 ps=19.29 w=19 l=1
X660 AVOUT1.t14 a_2308_n4916.t5 VSS.t127 sky130_fd_pr__res_high_po_0p69 l=12.22
X661 a_n2121_10269# a_n2577_9801# VDD.t46 VDD.t45 sky130_fd_pr__pfet_g5v0d10v5 ad=0.2142 pd=1.99 as=0.2142 ps=1.99 w=0.42 l=1
X662 x6.V1.t36 x9.V2.t23 VSS.t114 sky130_fd_pr__res_high_po_0p69 l=12.22
X663 x3.R1.t1 x8.V2.t1 VSS.t6 sky130_fd_pr__res_high_po_0p69 l=12.22
X664 AVOUT1.t29 a_6164_n4916.t26 VSS.t210 sky130_fd_pr__res_high_po_0p69 l=12.22
X665 a_n2577_n183# a_n2603_n130# DVSS.t183 DVSS.t182 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X666 x5.V2.t57 x4.V2.t58 VSS.t57 sky130_fd_pr__res_high_po_0p69 l=12.22
X667 x6.V1.t4 D93v3.t28 a_16261_n9984.t14 VSS.t21 sky130_fd_pr__nfet_g5v0d10v5 ad=0.638 pd=4.69 as=0.638 ps=4.69 w=4.4 l=1
X668 a_862_n3536# D03v3.t3 x4.V2.t59 VSS.t146 sky130_fd_pr__nfet_g5v0d10v5 ad=1.3833 pd=10.12 as=1.3833 ps=10.12 w=4.77 l=1
X669 ia_opamp_0.V2.t25 a_11509_n9984# VSS.t192 sky130_fd_pr__res_high_po_0p69 l=12.22
X670 a_7399_764.t3 V1.t0 a_6863_764.t1 VSS.t171 sky130_fd_pr__nfet_g5v0d10v5 ad=4.785 pd=33.58 as=4.785 ps=33.58 w=16.5 l=1
X671 DVSS.t246 a_n2559_n4073# a_n2121_n4707# DVSS.t245 sky130_fd_pr__nfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.21 ps=1.78 w=1.5 l=0.5
X672 x3.R1.t44 x8.V2.t42 VSS.t29 sky130_fd_pr__res_high_po_0p69 l=12.22
X673 x5.V2.t65 x4.V2.t66 VSS.t157 sky130_fd_pr__res_high_po_0p69 l=12.22
X674 x3.R1.t66 D93v3.t29 a_16261_n4916.t23 VSS.t21 sky130_fd_pr__nfet_g5v0d10v5 ad=0.638 pd=4.69 as=0.638 ps=4.69 w=4.4 l=1
X675 VOUT.t23 a_11509_n4916# VSS.t192 sky130_fd_pr__res_high_po_0p69 l=12.22
X676 a_n1825_4654# a_n2121_5277# VDD.t195 VDD.t102 sky130_fd_pr__pfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.24375 ps=1.825 w=1.5 l=0.5
X677 VDD.t166 a_n1825_n2834# D63v3.t1 VDD.t88 sky130_fd_pr__pfet_g5v0d10v5 ad=0.24375 pd=1.825 as=0.3975 ps=3.53 w=1.5 l=0.5
X678 a_3720_n9984.t3 D33v3.t16 x5.V2.t18 VSS.t89 sky130_fd_pr__nfet_g5v0d10v5 ad=0.6351 pd=4.67 as=0.6351 ps=4.67 w=4.38 l=1
X679 DVSS.t97 a_n2559_n6569# a_n2603_n7618# DVSS.t96 sky130_fd_pr__nfet_01v8 ad=0.1176 pd=1.12 as=0.2478 ps=2.27 w=0.84 l=0.15
X680 ia_opamp_0.V2.t22 a_16261_n9984.t12 VSS.t198 sky130_fd_pr__res_high_po_0p69 l=12.22
X681 a_3720_n4916.t2 D33v3.t17 x4.V2.t19 VSS.t89 sky130_fd_pr__nfet_g5v0d10v5 ad=0.6351 pd=4.67 as=0.6351 ps=4.67 w=4.38 l=1
X682 x8.V2.t46 a_10583_764.t7 VDD.t150 VDD.t149 sky130_fd_pr__pfet_g5v0d10v5 ad=2.755 pd=19.29 as=2.755 ps=19.29 w=19 l=1
X683 VOUT.t25 a_16261_n4916.t12 VSS.t198 sky130_fd_pr__res_high_po_0p69 l=12.22
X684 x3.R1.t23 x8.V2.t19 VSS.t118 sky130_fd_pr__res_high_po_0p69 l=12.22
X685 VDD.t216 DVSS.t314 VDD.t215 VDD.t214 sky130_fd_pr__pfet_g5v0d10v5 ad=0.265 pd=2.53 as=0 ps=0 w=1 l=1
X686 DVSS.t35 D5.t1 sky130_fd_pr__diode_pw2nd_11v0 perim=3.16e+06 area=6.072e+11
X687 x5.V2.t63 x4.V2.t64 VSS.t199 sky130_fd_pr__res_high_po_0p69 l=12.22
X688 x3.R1.t48 x8.V2.t48 VSS.t51 sky130_fd_pr__res_high_po_0p69 l=12.22
X689 ia_opamp_0.V2.t3 a_16261_n9984.t3 VSS.t36 sky130_fd_pr__res_high_po_0p69 l=12.22
X690 AVOUT1.t7 a_4215_764.t7 VDD.t22 VDD.t21 sky130_fd_pr__pfet_g5v0d10v5 ad=2.755 pd=19.29 as=5.51 ps=38.58 w=19 l=1
X691 x5.V2.t20 x4.V2.t21 VSS.t107 sky130_fd_pr__res_high_po_0p69 l=12.22
X692 VDD.t219 DVSS.t315 VDD.t218 VDD.t217 sky130_fd_pr__pfet_g5v0d10v5 ad=0.265 pd=2.53 as=0 ps=0 w=1 l=1
X693 x5.V2.t64 x4.V2.t65 VSS.t43 sky130_fd_pr__res_high_po_0p69 l=12.22
X694 a_n2121_12765# a_n2577_12297# VDD.t201 VDD.t200 sky130_fd_pr__pfet_g5v0d10v5 ad=0.2142 pd=1.99 as=0.2142 ps=1.99 w=0.42 l=1
X695 x3.R1.t61 x8.V2.t56 VSS.t94 sky130_fd_pr__res_high_po_0p69 l=12.22
X696 VOUT.t24 a_16261_n4916.t11 VSS.t36 sky130_fd_pr__res_high_po_0p69 l=12.22
X697 x6.V1.t35 x9.V2.t22 VSS.t6 sky130_fd_pr__res_high_po_0p69 l=12.22
X698 a_6598_281.t0 AVOUT2.t27 VSS.t224 sky130_fd_pr__res_high_po_0p69 l=3.2
X699 x6.V1.t37 x9.V2.t24 VSS.t29 sky130_fd_pr__res_high_po_0p69 l=12.22
X700 x3.R1.t7 x8.V2.t7 VSS.t8 sky130_fd_pr__res_high_po_0p69 l=12.22
X701 x3.R1.t2 x8.V2.t2 VSS.t7 sky130_fd_pr__res_high_po_0p69 l=12.22
X702 a_6164_n9984.t5 D43v3.t26 x5.V2.t10 VSS.t55 sky130_fd_pr__nfet_g5v0d10v5 ad=0.638 pd=4.69 as=0.638 ps=4.69 w=4.4 l=1
X703 amp_biases_0.ibias3.t1 amp_biases_0.ibias3.t0 VSS.t17 VSS.t16 sky130_fd_pr__nfet_g5v0d10v5 ad=4.4776 pd=31.46 as=4.4776 ps=31.46 w=15.44 l=1
X704 x3.R1.t35 x8.V2.t31 VSS.t170 sky130_fd_pr__res_high_po_0p69 l=12.22
X705 x5.V2.t70 x4.V2.t71 VSS.t141 sky130_fd_pr__res_high_po_0p69 l=12.22
X706 DVSS.t113 a_n1825_14638# sky130_fd_sc_hvl__lsbuflv2hv_1_0[10].X.t0 DVSS.t112 sky130_fd_pr__nfet_g5v0d10v5 ad=0.121875 pd=1.075 as=0.19875 ps=2.03 w=0.75 l=0.5
X707 a_13817_n9984.t12 D83v3.t10 x6.V1.t76 VSS.t233 sky130_fd_pr__nfet_g5v0d10v5 ad=1.2702 pd=9.34 as=0.6351 ps=4.67 w=4.38 l=1
X708 a_6164_n4916.t6 D43v3.t27 x4.V2.t22 VSS.t55 sky130_fd_pr__nfet_g5v0d10v5 ad=0.638 pd=4.69 as=0.638 ps=4.69 w=4.4 l=1
X709 x5.V2.t7 x4.V2.t8 VSS.t38 sky130_fd_pr__res_high_po_0p69 l=12.22
X710 a_10583_764.t1 a_9789_764.t6 VDD.t67 VDD.t66 sky130_fd_pr__pfet_g5v0d10v5 ad=2.175 pd=15.29 as=4.35 ps=30.58 w=15 l=1
X711 x6.V1.t43 x9.V2.t30 VSS.t118 sky130_fd_pr__res_high_po_0p69 l=12.22
X712 a_13817_n4916.t11 D83v3.t11 x3.R1.t63 VSS.t233 sky130_fd_pr__nfet_g5v0d10v5 ad=1.2702 pd=9.34 as=0.6351 ps=4.67 w=4.38 l=1
X713 AVOUT2.t4 a_7399_764.t6 VDD.t26 VDD.t25 sky130_fd_pr__pfet_g5v0d10v5 ad=2.755 pd=19.29 as=2.755 ps=19.29 w=19 l=1
X714 DVSS.t161 a_n2559_n9065# a_n2121_n9699# DVSS.t160 sky130_fd_pr__nfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.21 ps=1.78 w=1.5 l=0.5
X715 DVSS.t159 a_n2559_n9065# a_n2121_n9699# DVSS.t158 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.3975 ps=3.53 w=1.5 l=0.5
X716 x6.V1.t13 x9.V2.t7 VSS.t51 sky130_fd_pr__res_high_po_0p69 l=12.22
X717 AVOUT2.t3 a_6164_n9984.t1 VSS.t46 sky130_fd_pr__res_high_po_0p69 l=12.22
X718 a_n2577_7305# a_n2603_7358# DVSS.t231 DVSS.t229 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X719 x6.V1.t20 x9.V2.t10 VSS.t94 sky130_fd_pr__res_high_po_0p69 l=12.22
X720 AVOUT1.t25 a_6164_n4916.t23 VSS.t46 sky130_fd_pr__res_high_po_0p69 l=12.22
X721 AVOUT2.t2 a_3720_n9984.t1 VSS.t45 sky130_fd_pr__res_high_po_0p69 l=12.22
X722 VDD.t170 a_13767_764.t7 x9.V2.t50 VDD.t169 sky130_fd_pr__pfet_g5v0d10v5 ad=5.51 pd=38.58 as=2.755 ps=19.29 w=19 l=1
X723 x6.V1.t1 x9.V2.t0 VSS.t8 sky130_fd_pr__res_high_po_0p69 l=12.22
X724 AVOUT2.t17 a_6164_n9984.t20 VSS.t9 sky130_fd_pr__res_high_po_0p69 l=12.22
X725 x5.V2.t4 x4.V2.t4 VSS.t14 sky130_fd_pr__res_high_po_0p69 l=12.22
X726 a_n2559_5911# D3.t2 DVDD.t17 DVDD.t16 sky130_fd_pr__pfet_01v8_hvt ad=0.2478 pd=2.27 as=0.1176 ps=1.12 w=0.84 l=0.15
X727 DVSS.t216 a_n2559_13399# a_n2121_12765# DVSS.t215 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X728 a_n2559_919# D5.t2 DVDD.t5 DVDD.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.2478 pd=2.27 as=0.1176 ps=1.12 w=0.84 l=0.15
X729 AVOUT1.t9 a_3720_n4916.t1 VSS.t45 sky130_fd_pr__res_high_po_0p69 l=12.22
X730 x6.V1.t12 x9.V2.t6 VSS.t7 sky130_fd_pr__res_high_po_0p69 l=12.22
X731 AVOUT1.t0 a_6164_n4916.t0 VSS.t9 sky130_fd_pr__res_high_po_0p69 l=12.22
X732 VDD.t28 a_7399_764.t7 AVOUT2.t5 VDD.t27 sky130_fd_pr__pfet_g5v0d10v5 ad=2.755 pd=19.29 as=2.755 ps=19.29 w=19 l=1
X733 x6.V1.t63 x9.V2.t44 VSS.t170 sky130_fd_pr__res_high_po_0p69 l=12.22
X734 DVSS.t177 a_n2603_4862# a_n2577_4809# DVSS.t176 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X735 a_n1825_n338# a_n2121_285# DVSS.t53 DVSS.t52 sky130_fd_pr__nfet_g5v0d10v5 ad=0.19875 pd=2.03 as=0.121875 ps=1.075 w=0.75 l=0.5
X736 a_n2577_9801# a_n2603_9854# DVSS.t147 DVSS.t146 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X737 x3.R1.t4 x8.V2.t4 VSS.t39 sky130_fd_pr__res_high_po_0p69 l=12.22
X738 DVSS.t171 a_n2603_14846# a_n2577_14793# DVSS.t170 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X739 a_2622_12748.t2 a_2622_12748.t1 VSS.t216 VSS.t215 sky130_fd_pr__nfet_g5v0d10v5 ad=2.2388 pd=15.73 as=2.2388 ps=15.73 w=15.44 l=1
X740 ia_opamp_0.V2.t10 a_13817_n9984.t0 VSS.t10 sky130_fd_pr__res_high_po_0p69 l=12.22
X741 x5.V2.t21 D43v3.t28 a_6164_n9984.t4 VSS.t108 sky130_fd_pr__nfet_g5v0d10v5 ad=0.638 pd=4.69 as=0.638 ps=4.69 w=4.4 l=1
X742 DVSS.t95 a_n2559_n6569# a_n2121_n7203# DVSS.t94 sky130_fd_pr__nfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.21 ps=1.78 w=1.5 l=0.5
X743 amp_biases_0.ibias5.t2 a_204_12823.t15 VDD.t185 VDD.t184 sky130_fd_pr__pfet_g5v0d10v5 ad=2.175 pd=15.29 as=2.175 ps=15.29 w=15 l=1
X744 x4.V2.t23 D43v3.t29 a_6164_n4916.t5 VSS.t108 sky130_fd_pr__nfet_g5v0d10v5 ad=0.638 pd=4.69 as=0.638 ps=4.69 w=4.4 l=1
X745 VOUT.t0 a_13817_n4916.t0 VSS.t10 sky130_fd_pr__res_high_po_0p69 l=12.22
X746 a_n1825_7150# a_n2121_7773# VDD.t151 VDD.t41 sky130_fd_pr__pfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.24375 ps=1.825 w=1.5 l=0.5
X747 DVSS.t193 a_n1825_n2834# D63v3.t0 DVSS.t192 sky130_fd_pr__nfet_g5v0d10v5 ad=0.121875 pd=1.075 as=0.19875 ps=2.03 w=0.75 l=0.5
X748 x6.V1.t74 D83v3.t12 a_13817_n9984.t10 VSS.t231 sky130_fd_pr__nfet_g5v0d10v5 ad=0.6351 pd=4.67 as=0.6351 ps=4.67 w=4.38 l=1
X749 x5.V2.t33 x4.V2.t32 VSS.t145 sky130_fd_pr__res_high_po_0p69 l=12.22
X750 DVSS.t157 a_n2559_n9065# a_n2603_n10114# DVSS.t156 sky130_fd_pr__nfet_01v8 ad=0.1176 pd=1.12 as=0.2478 ps=2.27 w=0.84 l=0.15
X751 ia_opamp_0.V2.t24 a_13817_n9984.t8 VSS.t225 sky130_fd_pr__res_high_po_0p69 l=12.22
X752 x3.R1.t60 D83v3.t13 a_13817_n4916.t9 VSS.t231 sky130_fd_pr__nfet_g5v0d10v5 ad=0.6351 pd=4.67 as=0.6351 ps=4.67 w=4.38 l=1
X753 DVSS.t119 a_n2559_15895# a_n2121_15261# DVSS.t118 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X754 a_n2559_3415# D4.t2 DVDD.t21 DVDD.t20 sky130_fd_pr__pfet_01v8_hvt ad=0.2478 pd=2.27 as=0.1176 ps=1.12 w=0.84 l=0.15
X755 x3.R1.t57 x8.V2.t55 VSS.t178 sky130_fd_pr__res_high_po_0p69 l=12.22
X756 x6.V1.t75 D83v3.t14 a_13817_n9984.t11 VSS.t229 sky130_fd_pr__nfet_g5v0d10v5 ad=0.6351 pd=4.67 as=0.6351 ps=4.67 w=4.38 l=1
X757 VOUT.t28 a_13817_n4916.t6 VSS.t225 sky130_fd_pr__res_high_po_0p69 l=12.22
X758 a_n2121_15261# a_n2559_15895# DVSS.t115 DVSS.t114 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X759 DVSS.t274 VDD.t248 DVSS.t273 DVSS.t272 sky130_fd_pr__nfet_g5v0d10v5 ad=0.19875 pd=2.03 as=0 ps=0 w=0.75 l=1
X760 VDD.t222 DVSS.t316 VDD.t221 VDD.t220 sky130_fd_pr__pfet_g5v0d10v5 ad=0.265 pd=2.53 as=0 ps=0 w=1 l=1
X761 DVSS.t230 a_n2603_7358# a_n2577_7305# DVSS.t229 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X762 AVOUT2.t28 a_2308_n9984.t6 VSS.t226 sky130_fd_pr__res_high_po_0p69 l=12.22
X763 VDD.t106 DVSS.t317 VDD.t105 VDD.t104 sky130_fd_pr__pfet_g5v0d10v5 ad=0.265 pd=2.53 as=0 ps=0 w=1 l=1
X764 x3.R1.t43 x8.V2.t41 VSS.t137 sky130_fd_pr__res_high_po_0p69 l=12.22
X765 VDD.t187 a_204_12823.t16 amp_biases_0.ibias4.t2 VDD.t186 sky130_fd_pr__pfet_g5v0d10v5 ad=2.175 pd=15.29 as=2.175 ps=15.29 w=15 l=1
X766 x3.R1.t58 D83v3.t15 a_13817_n4916.t7 VSS.t229 sky130_fd_pr__nfet_g5v0d10v5 ad=0.6351 pd=4.67 as=0.6351 ps=4.67 w=4.38 l=1
X767 a_n2121_15261# a_n2577_14793# VDD.t95 VDD.t94 sky130_fd_pr__pfet_g5v0d10v5 ad=0.2142 pd=1.99 as=0.2142 ps=1.99 w=0.42 l=1
X768 x6.V1.t66 x9.V2.t48 VSS.t39 sky130_fd_pr__res_high_po_0p69 l=12.22
X769 AVOUT1.t31 a_2308_n4916.t6 VSS.t226 sky130_fd_pr__res_high_po_0p69 l=12.22
X770 a_230_281.t1 a_1031_764.t2 sky130_fd_pr__cap_mim_m3_1 l=6.9 w=6.9
X771 x5.V2.t66 x4.V2.t67 VSS.t85 sky130_fd_pr__res_high_po_0p69 l=12.22
X772 amp_biases_0.ibias4.t1 amp_biases_0.ibias4.t0 VSS.t176 VSS.t175 sky130_fd_pr__nfet_g5v0d10v5 ad=4.4776 pd=31.46 as=4.4776 ps=31.46 w=15.44 l=1
X773 DVSS.t127 a_n2603_n5122# a_n2577_n5175# DVSS.t126 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X774 a_13767_764.t0 a_12973_764.t6 VDD.t52 VDD.t51 sky130_fd_pr__pfet_g5v0d10v5 ad=2.175 pd=15.29 as=4.35 ps=30.58 w=15 l=1
X775 a_n1825_9646# a_n2121_10269# VDD.t126 VDD.t31 sky130_fd_pr__pfet_g5v0d10v5 ad=0.3975 pd=3.53 as=0.24375 ps=1.825 w=1.5 l=0.5
X776 VDD.t1 a_n1825_n10322# D93v3.t1 VDD.t0 sky130_fd_pr__pfet_g5v0d10v5 ad=0.24375 pd=1.825 as=0.3975 ps=3.53 w=1.5 l=0.5
X777 a_n2121_2781# a_n2559_3415# DVSS.t204 DVSS.t203 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X778 VSS.t238 a_2622_12748.t3 a_2564_12836# VSS.t237 sky130_fd_pr__nfet_g5v0d10v5 ad=2.2388 pd=15.73 as=2.2388 ps=15.73 w=15.44 l=1
X779 x6.V1.t68 x9.V2.t52 VSS.t178 sky130_fd_pr__res_high_po_0p69 l=12.22
X780 DVSS.t21 D8.t2 sky130_fd_pr__diode_pw2nd_11v0 perim=3.16e+06 area=6.072e+11
X781 x3.R1.t54 x8.V2.t54 VSS.t160 sky130_fd_pr__res_high_po_0p69 l=12.22
X782 ia_opamp_0.V2.t26 a_12405_n9984.t6 VSS.t15 sky130_fd_pr__res_high_po_0p69 l=12.22
X783 a_n2577_n2679# a_n2603_n2626# DVSS.t139 DVSS.t138 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X784 x6.V1.t67 x9.V2.t51 VSS.t137 sky130_fd_pr__res_high_po_0p69 l=12.22
X785 x3.R1.t53 x8.V2.t53 VSS.t199 sky130_fd_pr__res_high_po_0p69 l=12.22
X786 ia_opamp_0.V2.t7 a_16261_n9984.t6 VSS.t95 sky130_fd_pr__res_high_po_0p69 l=12.22
X787 VOUT.t1 a_12405_n4916.t0 VSS.t15 sky130_fd_pr__res_high_po_0p69 l=12.22
X788 a_13817_n9984.t9 D83v3.t16 x6.V1.t73 VSS.t230 sky130_fd_pr__nfet_g5v0d10v5 ad=0.6351 pd=4.67 as=0.6351 ps=4.67 w=4.38 l=1
X789 VOUT.t7 a_16261_n4916.t2 VSS.t95 sky130_fd_pr__res_high_po_0p69 l=12.22
X790 VDD.t83 a_16951_764.t7 VOUT.t30 VDD.t82 sky130_fd_pr__pfet_g5v0d10v5 ad=5.51 pd=38.58 as=2.755 ps=19.29 w=19 l=1
X791 VDD.t227 a_1031_764.t7 ia_opamp_0.V2.t34 VDD.t226 sky130_fd_pr__pfet_g5v0d10v5 ad=5.51 pd=38.58 as=2.755 ps=19.29 w=19 l=1
X792 DVDD.t1 a_n2559_10903# a_n2603_9854# DVDD.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.12 as=0.2478 ps=2.27 w=0.84 l=0.15
X793 a_n2559_8407# D2.t2 DVDD.t11 DVDD.t10 sky130_fd_pr__pfet_01v8_hvt ad=0.2478 pd=2.27 as=0.1176 ps=1.12 w=0.84 l=0.15
X794 a_13817_n4916.t8 D83v3.t17 x3.R1.t59 VSS.t230 sky130_fd_pr__nfet_g5v0d10v5 ad=0.6351 pd=4.67 as=0.6351 ps=4.67 w=4.38 l=1
X795 x3.R1.t33 x8.V2.t28 VSS.t0 sky130_fd_pr__res_high_po_0p69 l=12.22
X796 x3.R1.t31 x8.V2.t26 VSS.t158 sky130_fd_pr__res_high_po_0p69 l=12.22
X797 x5.V2.t13 x4.V2.t14 VSS.t42 sky130_fd_pr__res_high_po_0p69 l=12.22
X798 a_n1825_2158# a_n2121_2781# DVSS.t195 DVSS.t194 sky130_fd_pr__nfet_g5v0d10v5 ad=0.19875 pd=2.03 as=0.121875 ps=1.075 w=0.75 l=0.5
X799 a_n2559_n1577# D6.t2 DVDD.t27 DVDD.t26 sky130_fd_pr__pfet_01v8_hvt ad=0.2478 pd=2.27 as=0.1176 ps=1.12 w=0.84 l=0.15
X800 x3.R1.t28 x8.V2.t23 VSS.t107 sky130_fd_pr__res_high_po_0p69 l=12.22
R0 x6.V1.n0 x6.V1.t94 491.978
R1 x6.V1.n158 x6.V1.t29 22.474
R2 x6.V1.n131 x6.V1.n129 20.8462
R3 x6.V1.n1 x6.V1.t81 20.705
R4 x6.V1.n3 x6.V1.t79 20.705
R5 x6.V1.n4 x6.V1.t13 20.705
R6 x6.V1.n5 x6.V1.t37 20.705
R7 x6.V1.n6 x6.V1.t10 20.705
R8 x6.V1.n7 x6.V1.t44 20.705
R9 x6.V1.n8 x6.V1.t38 20.705
R10 x6.V1.n9 x6.V1.t64 20.705
R11 x6.V1.n10 x6.V1.t8 20.705
R12 x6.V1.n11 x6.V1.t28 20.705
R13 x6.V1.n12 x6.V1.t89 20.705
R14 x6.V1.n13 x6.V1.t72 20.705
R15 x6.V1.n14 x6.V1.t66 20.705
R16 x6.V1.n15 x6.V1.t21 20.705
R17 x6.V1.n16 x6.V1.t31 20.705
R18 x6.V1.n17 x6.V1.t46 20.705
R19 x6.V1.n18 x6.V1.t88 20.705
R20 x6.V1.n19 x6.V1.t80 20.705
R21 x6.V1.n20 x6.V1.t40 20.705
R22 x6.V1.n21 x6.V1.t43 20.705
R23 x6.V1.n22 x6.V1.t35 20.705
R24 x6.V1.n23 x6.V1.t26 20.705
R25 x6.V1.n24 x6.V1.t52 20.705
R26 x6.V1.n25 x6.V1.t54 20.705
R27 x6.V1.n26 x6.V1.t50 20.705
R28 x6.V1.n27 x6.V1.t57 20.705
R29 x6.V1.n28 x6.V1.t34 20.705
R30 x6.V1.n29 x6.V1.t33 20.705
R31 x6.V1.n31 x6.V1.t49 20.705
R32 x6.V1.n32 x6.V1.t39 20.705
R33 x6.V1.n33 x6.V1.t90 20.705
R34 x6.V1.n34 x6.V1.t7 20.705
R35 x6.V1.n35 x6.V1.t93 20.705
R36 x6.V1.n36 x6.V1.t42 20.705
R37 x6.V1.n37 x6.V1.t16 20.705
R38 x6.V1.n38 x6.V1.t48 20.705
R39 x6.V1.n39 x6.V1.t67 20.705
R40 x6.V1.n40 x6.V1.t36 20.705
R41 x6.V1.n41 x6.V1.t92 20.705
R42 x6.V1.n42 x6.V1.t65 20.705
R43 x6.V1.n43 x6.V1.t87 20.705
R44 x6.V1.n44 x6.V1.t91 20.705
R45 x6.V1.n45 x6.V1.t78 20.705
R46 x6.V1.n46 x6.V1.t32 20.705
R47 x6.V1.n47 x6.V1.t20 20.705
R48 x6.V1.n48 x6.V1.t47 20.705
R49 x6.V1.n49 x6.V1.t12 20.705
R50 x6.V1.n50 x6.V1.t56 20.705
R51 x6.V1.n51 x6.V1.t30 20.705
R52 x6.V1.n52 x6.V1.t86 20.705
R53 x6.V1.n53 x6.V1.t62 20.705
R54 x6.V1.n54 x6.V1.t85 20.705
R55 x6.V1.n55 x6.V1.t24 20.705
R56 x6.V1.n56 x6.V1.t68 20.705
R57 x6.V1.n57 x6.V1.t19 20.705
R58 x6.V1.n58 x6.V1.t51 20.705
R59 x6.V1.n59 x6.V1.t9 20.705
R60 x6.V1.n60 x6.V1.t11 20.705
R61 x6.V1.n61 x6.V1.t84 20.705
R62 x6.V1.n62 x6.V1.t41 20.705
R63 x6.V1.n123 x6.V1.t63 20.705
R64 x6.V1.n124 x6.V1.t25 20.705
R65 x6.V1.n126 x6.V1.t45 20.705
R66 x6.V1.n30 x6.V1.t1 20.705
R67 x6.V1.n155 x6.V1.n154 19.9925
R68 x6.V1.n153 x6.V1.n152 19.9925
R69 x6.V1.n143 x6.V1.n142 19.9842
R70 x6.V1.n141 x6.V1.n140 19.9842
R71 x6.V1.n139 x6.V1.n138 19.9842
R72 x6.V1.n137 x6.V1.n136 19.9842
R73 x6.V1.n135 x6.V1.n134 19.9842
R74 x6.V1.n133 x6.V1.n132 19.9842
R75 x6.V1.n131 x6.V1.n130 19.9842
R76 x6.V1.n151 x6.V1.n150 19.9788
R77 x6.V1.n149 x6.V1.n148 19.9788
R78 x6.V1.n147 x6.V1.n146 19.9788
R79 x6.V1.n145 x6.V1.n144 19.9788
R80 x6.V1.n157 x6.V1.n156 19.0358
R81 x6.V1.n159 x6.V1.t53 17.8929
R82 x6.V1.n129 x6.V1.n128 15.5786
R83 x6.V1.n129 x6.V1.n0 7.09738
R84 x6.V1.n159 x6.V1.n158 5.42932
R85 x6.V1.n150 x6.V1.t73 3.77447
R86 x6.V1.n150 x6.V1.t59 3.77447
R87 x6.V1.n148 x6.V1.t60 3.77447
R88 x6.V1.n148 x6.V1.t75 3.77447
R89 x6.V1.n146 x6.V1.t77 3.77447
R90 x6.V1.n146 x6.V1.t58 3.77447
R91 x6.V1.n144 x6.V1.t76 3.77447
R92 x6.V1.n144 x6.V1.t74 3.77447
R93 x6.V1.n142 x6.V1.t55 3.75732
R94 x6.V1.n142 x6.V1.t3 3.75732
R95 x6.V1.n140 x6.V1.t0 3.75732
R96 x6.V1.n140 x6.V1.t22 3.75732
R97 x6.V1.n138 x6.V1.t71 3.75732
R98 x6.V1.n138 x6.V1.t4 3.75732
R99 x6.V1.n136 x6.V1.t6 3.75732
R100 x6.V1.n136 x6.V1.t70 3.75732
R101 x6.V1.n134 x6.V1.t23 3.75732
R102 x6.V1.n134 x6.V1.t5 3.75732
R103 x6.V1.n132 x6.V1.t61 3.75732
R104 x6.V1.n132 x6.V1.t18 3.75732
R105 x6.V1.n130 x6.V1.t2 3.75732
R106 x6.V1.n130 x6.V1.t27 3.75732
R107 x6.V1.n154 x6.V1.t17 3.55534
R108 x6.V1.n154 x6.V1.t83 3.55534
R109 x6.V1.n152 x6.V1.t15 3.55534
R110 x6.V1.n152 x6.V1.t14 3.55534
R111 x6.V1.n156 x6.V1.t82 3.39475
R112 x6.V1.n156 x6.V1.t69 3.39475
R113 x6.V1.n145 x6.V1.n143 1.55606
R114 x6.V1.n153 x6.V1.n151 1.55606
R115 x6.V1.n157 x6.V1.n155 1.55606
R116 x6.V1.n158 x6.V1.n157 1.55606
R117 x6.V1.n0 x6.V1 0.929667
R118 x6.V1.n147 x6.V1.n145 0.898069
R119 x6.V1.n151 x6.V1.n149 0.898069
R120 x6.V1.n133 x6.V1.n131 0.896333
R121 x6.V1.n135 x6.V1.n133 0.896333
R122 x6.V1.n137 x6.V1.n135 0.896333
R123 x6.V1.n139 x6.V1.n137 0.896333
R124 x6.V1.n143 x6.V1.n141 0.896333
R125 x6.V1.n155 x6.V1.n153 0.896333
R126 x6.V1.n141 x6.V1.n139 0.894597
R127 x6.V1.n149 x6.V1.n147 0.894597
R128 x6.V1.n63 x6.V1.n3 0.844944
R129 x6.V1.n128 x6.V1.n1 0.794713
R130 x6.V1.n63 x6.V1.n4 0.777392
R131 x6.V1.n64 x6.V1.n5 0.777392
R132 x6.V1.n65 x6.V1.n6 0.777392
R133 x6.V1.n66 x6.V1.n7 0.777392
R134 x6.V1.n67 x6.V1.n8 0.777392
R135 x6.V1.n68 x6.V1.n9 0.777392
R136 x6.V1.n69 x6.V1.n10 0.777392
R137 x6.V1.n70 x6.V1.n11 0.777392
R138 x6.V1.n71 x6.V1.n12 0.777392
R139 x6.V1.n72 x6.V1.n13 0.777392
R140 x6.V1.n73 x6.V1.n14 0.777392
R141 x6.V1.n74 x6.V1.n15 0.777392
R142 x6.V1.n75 x6.V1.n16 0.777392
R143 x6.V1.n76 x6.V1.n17 0.777392
R144 x6.V1.n77 x6.V1.n18 0.777392
R145 x6.V1.n78 x6.V1.n19 0.777392
R146 x6.V1.n79 x6.V1.n20 0.777392
R147 x6.V1.n80 x6.V1.n21 0.777392
R148 x6.V1.n81 x6.V1.n22 0.777392
R149 x6.V1.n82 x6.V1.n23 0.777392
R150 x6.V1.n83 x6.V1.n24 0.777392
R151 x6.V1.n84 x6.V1.n25 0.777392
R152 x6.V1.n85 x6.V1.n26 0.777392
R153 x6.V1.n86 x6.V1.n27 0.777392
R154 x6.V1.n87 x6.V1.n28 0.777392
R155 x6.V1.n88 x6.V1.n29 0.777392
R156 x6.V1.n90 x6.V1.n31 0.777392
R157 x6.V1.n91 x6.V1.n32 0.777392
R158 x6.V1.n92 x6.V1.n33 0.777392
R159 x6.V1.n93 x6.V1.n34 0.777392
R160 x6.V1.n94 x6.V1.n35 0.777392
R161 x6.V1.n95 x6.V1.n36 0.777392
R162 x6.V1.n96 x6.V1.n37 0.777392
R163 x6.V1.n97 x6.V1.n38 0.777392
R164 x6.V1.n98 x6.V1.n39 0.777392
R165 x6.V1.n99 x6.V1.n40 0.777392
R166 x6.V1.n100 x6.V1.n41 0.777392
R167 x6.V1.n101 x6.V1.n42 0.777392
R168 x6.V1.n102 x6.V1.n43 0.777392
R169 x6.V1.n103 x6.V1.n44 0.777392
R170 x6.V1.n104 x6.V1.n45 0.777392
R171 x6.V1.n105 x6.V1.n46 0.777392
R172 x6.V1.n106 x6.V1.n47 0.777392
R173 x6.V1.n107 x6.V1.n48 0.777392
R174 x6.V1.n108 x6.V1.n49 0.777392
R175 x6.V1.n109 x6.V1.n50 0.777392
R176 x6.V1.n110 x6.V1.n51 0.777392
R177 x6.V1.n111 x6.V1.n52 0.777392
R178 x6.V1.n112 x6.V1.n53 0.777392
R179 x6.V1.n113 x6.V1.n54 0.777392
R180 x6.V1.n114 x6.V1.n55 0.777392
R181 x6.V1.n115 x6.V1.n56 0.777392
R182 x6.V1.n116 x6.V1.n57 0.777392
R183 x6.V1.n117 x6.V1.n58 0.777392
R184 x6.V1.n118 x6.V1.n59 0.777392
R185 x6.V1.n119 x6.V1.n60 0.777392
R186 x6.V1.n120 x6.V1.n61 0.777392
R187 x6.V1.n121 x6.V1.n62 0.777392
R188 x6.V1.n123 x6.V1.n122 0.777392
R189 x6.V1.n124 x6.V1.n2 0.777392
R190 x6.V1.n127 x6.V1.n126 0.777392
R191 x6.V1.n89 x6.V1.n30 0.777392
R192 x6.V1.n125 x6.V1.n3 0.74147
R193 x6.V1.n125 x6.V1.n4 0.74147
R194 x6.V1.n125 x6.V1.n5 0.74147
R195 x6.V1.n125 x6.V1.n6 0.74147
R196 x6.V1.n125 x6.V1.n7 0.74147
R197 x6.V1.n125 x6.V1.n8 0.74147
R198 x6.V1.n125 x6.V1.n9 0.74147
R199 x6.V1.n125 x6.V1.n10 0.74147
R200 x6.V1.n125 x6.V1.n11 0.74147
R201 x6.V1.n125 x6.V1.n12 0.74147
R202 x6.V1.n125 x6.V1.n13 0.74147
R203 x6.V1.n125 x6.V1.n14 0.74147
R204 x6.V1.n125 x6.V1.n15 0.74147
R205 x6.V1.n125 x6.V1.n16 0.74147
R206 x6.V1.n125 x6.V1.n17 0.74147
R207 x6.V1.n125 x6.V1.n18 0.74147
R208 x6.V1.n125 x6.V1.n19 0.74147
R209 x6.V1.n125 x6.V1.n20 0.74147
R210 x6.V1.n125 x6.V1.n21 0.74147
R211 x6.V1.n125 x6.V1.n22 0.74147
R212 x6.V1.n125 x6.V1.n23 0.74147
R213 x6.V1.n125 x6.V1.n24 0.74147
R214 x6.V1.n125 x6.V1.n25 0.74147
R215 x6.V1.n125 x6.V1.n26 0.74147
R216 x6.V1.n125 x6.V1.n27 0.74147
R217 x6.V1.n125 x6.V1.n28 0.74147
R218 x6.V1.n125 x6.V1.n29 0.74147
R219 x6.V1.n125 x6.V1.n30 0.74147
R220 x6.V1.n125 x6.V1.n31 0.74147
R221 x6.V1.n125 x6.V1.n32 0.74147
R222 x6.V1.n125 x6.V1.n33 0.74147
R223 x6.V1.n125 x6.V1.n34 0.74147
R224 x6.V1.n125 x6.V1.n35 0.74147
R225 x6.V1.n125 x6.V1.n36 0.74147
R226 x6.V1.n125 x6.V1.n37 0.74147
R227 x6.V1.n125 x6.V1.n38 0.74147
R228 x6.V1.n125 x6.V1.n39 0.74147
R229 x6.V1.n125 x6.V1.n40 0.74147
R230 x6.V1.n125 x6.V1.n41 0.74147
R231 x6.V1.n125 x6.V1.n42 0.74147
R232 x6.V1.n125 x6.V1.n43 0.74147
R233 x6.V1.n125 x6.V1.n44 0.74147
R234 x6.V1.n125 x6.V1.n45 0.74147
R235 x6.V1.n125 x6.V1.n46 0.74147
R236 x6.V1.n125 x6.V1.n47 0.74147
R237 x6.V1.n125 x6.V1.n48 0.74147
R238 x6.V1.n125 x6.V1.n49 0.74147
R239 x6.V1.n125 x6.V1.n50 0.74147
R240 x6.V1.n125 x6.V1.n51 0.74147
R241 x6.V1.n125 x6.V1.n52 0.74147
R242 x6.V1.n125 x6.V1.n53 0.74147
R243 x6.V1.n125 x6.V1.n54 0.74147
R244 x6.V1.n125 x6.V1.n55 0.74147
R245 x6.V1.n125 x6.V1.n56 0.74147
R246 x6.V1.n125 x6.V1.n57 0.74147
R247 x6.V1.n125 x6.V1.n58 0.74147
R248 x6.V1.n125 x6.V1.n59 0.74147
R249 x6.V1.n125 x6.V1.n60 0.74147
R250 x6.V1.n125 x6.V1.n61 0.74147
R251 x6.V1.n125 x6.V1.n62 0.74147
R252 x6.V1.n125 x6.V1.n123 0.74147
R253 x6.V1.n125 x6.V1.n124 0.74147
R254 x6.V1.n126 x6.V1.n125 0.74147
R255 x6.V1.n125 x6.V1.n1 0.74147
R256 x6.V1 x6.V1.n159 0.558313
R257 x6.V1.n127 x6.V1.n2 0.068052
R258 x6.V1.n122 x6.V1.n2 0.068052
R259 x6.V1.n122 x6.V1.n121 0.068052
R260 x6.V1.n121 x6.V1.n120 0.068052
R261 x6.V1.n120 x6.V1.n119 0.068052
R262 x6.V1.n119 x6.V1.n118 0.068052
R263 x6.V1.n118 x6.V1.n117 0.068052
R264 x6.V1.n117 x6.V1.n116 0.068052
R265 x6.V1.n116 x6.V1.n115 0.068052
R266 x6.V1.n115 x6.V1.n114 0.068052
R267 x6.V1.n114 x6.V1.n113 0.068052
R268 x6.V1.n113 x6.V1.n112 0.068052
R269 x6.V1.n112 x6.V1.n111 0.068052
R270 x6.V1.n111 x6.V1.n110 0.068052
R271 x6.V1.n110 x6.V1.n109 0.068052
R272 x6.V1.n109 x6.V1.n108 0.068052
R273 x6.V1.n108 x6.V1.n107 0.068052
R274 x6.V1.n107 x6.V1.n106 0.068052
R275 x6.V1.n106 x6.V1.n105 0.068052
R276 x6.V1.n105 x6.V1.n104 0.068052
R277 x6.V1.n104 x6.V1.n103 0.068052
R278 x6.V1.n103 x6.V1.n102 0.068052
R279 x6.V1.n102 x6.V1.n101 0.068052
R280 x6.V1.n101 x6.V1.n100 0.068052
R281 x6.V1.n100 x6.V1.n99 0.068052
R282 x6.V1.n99 x6.V1.n98 0.068052
R283 x6.V1.n98 x6.V1.n97 0.068052
R284 x6.V1.n97 x6.V1.n96 0.068052
R285 x6.V1.n96 x6.V1.n95 0.068052
R286 x6.V1.n95 x6.V1.n94 0.068052
R287 x6.V1.n94 x6.V1.n93 0.068052
R288 x6.V1.n93 x6.V1.n92 0.068052
R289 x6.V1.n92 x6.V1.n91 0.068052
R290 x6.V1.n91 x6.V1.n90 0.068052
R291 x6.V1.n90 x6.V1.n89 0.068052
R292 x6.V1.n89 x6.V1.n88 0.068052
R293 x6.V1.n88 x6.V1.n87 0.068052
R294 x6.V1.n87 x6.V1.n86 0.068052
R295 x6.V1.n86 x6.V1.n85 0.068052
R296 x6.V1.n85 x6.V1.n84 0.068052
R297 x6.V1.n84 x6.V1.n83 0.068052
R298 x6.V1.n83 x6.V1.n82 0.068052
R299 x6.V1.n82 x6.V1.n81 0.068052
R300 x6.V1.n81 x6.V1.n80 0.068052
R301 x6.V1.n80 x6.V1.n79 0.068052
R302 x6.V1.n79 x6.V1.n78 0.068052
R303 x6.V1.n78 x6.V1.n77 0.068052
R304 x6.V1.n77 x6.V1.n76 0.068052
R305 x6.V1.n76 x6.V1.n75 0.068052
R306 x6.V1.n75 x6.V1.n74 0.068052
R307 x6.V1.n74 x6.V1.n73 0.068052
R308 x6.V1.n73 x6.V1.n72 0.068052
R309 x6.V1.n72 x6.V1.n71 0.068052
R310 x6.V1.n71 x6.V1.n70 0.068052
R311 x6.V1.n70 x6.V1.n69 0.068052
R312 x6.V1.n69 x6.V1.n68 0.068052
R313 x6.V1.n68 x6.V1.n67 0.068052
R314 x6.V1.n67 x6.V1.n66 0.068052
R315 x6.V1.n66 x6.V1.n65 0.068052
R316 x6.V1.n65 x6.V1.n64 0.068052
R317 x6.V1.n64 x6.V1.n63 0.068052
R318 x6.V1.n128 x6.V1.n127 0.0507309
R319 x9.V2.n137 x9.V2.t70 491.709
R320 x9.V2.n135 x9.V2.t17 39.1599
R321 x9.V2.n125 x9.V2.t59 20.7986
R322 x9.V2.n4 x9.V2.t57 20.7986
R323 x9.V2.n5 x9.V2.t7 20.7986
R324 x9.V2.n6 x9.V2.t24 20.7986
R325 x9.V2.n7 x9.V2.t4 20.7986
R326 x9.V2.n8 x9.V2.t31 20.7986
R327 x9.V2.n9 x9.V2.t25 20.7986
R328 x9.V2.n10 x9.V2.t46 20.7986
R329 x9.V2.n11 x9.V2.t2 20.7986
R330 x9.V2.n12 x9.V2.t15 20.7986
R331 x9.V2.n13 x9.V2.t65 20.7986
R332 x9.V2.n14 x9.V2.t53 20.7986
R333 x9.V2.n15 x9.V2.t48 20.7986
R334 x9.V2.n16 x9.V2.t11 20.7986
R335 x9.V2.n17 x9.V2.t18 20.7986
R336 x9.V2.n18 x9.V2.t33 20.7986
R337 x9.V2.n19 x9.V2.t64 20.7986
R338 x9.V2.n20 x9.V2.t58 20.7986
R339 x9.V2.n21 x9.V2.t27 20.7986
R340 x9.V2.n22 x9.V2.t30 20.7986
R341 x9.V2.n23 x9.V2.t22 20.7986
R342 x9.V2.n24 x9.V2.t14 20.7986
R343 x9.V2.n25 x9.V2.t39 20.7986
R344 x9.V2.n26 x9.V2.t40 20.7986
R345 x9.V2.n27 x9.V2.t37 20.7986
R346 x9.V2.n28 x9.V2.t42 20.7986
R347 x9.V2.n29 x9.V2.t21 20.7986
R348 x9.V2.n30 x9.V2.t20 20.7986
R349 x9.V2.n32 x9.V2.t36 20.7986
R350 x9.V2.n33 x9.V2.t26 20.7986
R351 x9.V2.n34 x9.V2.t66 20.7986
R352 x9.V2.n35 x9.V2.t1 20.7986
R353 x9.V2.n36 x9.V2.t69 20.7986
R354 x9.V2.n37 x9.V2.t29 20.7986
R355 x9.V2.n38 x9.V2.t8 20.7986
R356 x9.V2.n39 x9.V2.t35 20.7986
R357 x9.V2.n40 x9.V2.t51 20.7986
R358 x9.V2.n41 x9.V2.t23 20.7986
R359 x9.V2.n42 x9.V2.t68 20.7986
R360 x9.V2.n43 x9.V2.t47 20.7986
R361 x9.V2.n44 x9.V2.t63 20.7986
R362 x9.V2.n45 x9.V2.t67 20.7986
R363 x9.V2.n46 x9.V2.t56 20.7986
R364 x9.V2.n47 x9.V2.t19 20.7986
R365 x9.V2.n48 x9.V2.t10 20.7986
R366 x9.V2.n49 x9.V2.t34 20.7986
R367 x9.V2.n50 x9.V2.t6 20.7986
R368 x9.V2.n51 x9.V2.t41 20.7986
R369 x9.V2.n52 x9.V2.t16 20.7986
R370 x9.V2.n53 x9.V2.t62 20.7986
R371 x9.V2.n104 x9.V2.t43 20.7986
R372 x9.V2.n105 x9.V2.t61 20.7986
R373 x9.V2.n127 x9.V2.t12 20.7986
R374 x9.V2.n106 x9.V2.t52 20.7986
R375 x9.V2.n107 x9.V2.t9 20.7986
R376 x9.V2.n108 x9.V2.t38 20.7986
R377 x9.V2.n109 x9.V2.t3 20.7986
R378 x9.V2.n110 x9.V2.t5 20.7986
R379 x9.V2.n111 x9.V2.t60 20.7986
R380 x9.V2.n112 x9.V2.t28 20.7986
R381 x9.V2.n113 x9.V2.t44 20.7986
R382 x9.V2.n114 x9.V2.t13 20.7986
R383 x9.V2.n115 x9.V2.t32 20.7986
R384 x9.V2.n132 x9.V2.n131 10.6258
R385 x9.V2.n1 x9.V2.n0 10.6258
R386 x9.V2.n137 x9.V2.n136 6.89614
R387 x9.V2.n133 x9.V2.n1 6.47346
R388 x9.V2.n133 x9.V2.n132 6.27518
R389 x9.V2.n136 x9.V2.n135 6.23929
R390 x9.V2.n130 x9.V2.n1 5.09996
R391 x9.V2.n132 x9.V2.n130 4.87014
R392 x9.V2.n130 x9.V2.n129 4.64492
R393 x9.V2.n135 x9.V2.t45 4.35292
R394 x9.V2.n134 x9.V2 2.58592
R395 x9.V2.n131 x9.V2.t50 1.45813
R396 x9.V2.n131 x9.V2.t49 1.45813
R397 x9.V2.n0 x9.V2.t54 1.45813
R398 x9.V2.n0 x9.V2.t55 1.45813
R399 x9.V2.n125 x9.V2.n124 0.843052
R400 x9.V2.n54 x9.V2.n4 0.843052
R401 x9.V2.n124 x9.V2.n115 0.7755
R402 x9.V2.n123 x9.V2.n114 0.7755
R403 x9.V2.n122 x9.V2.n113 0.7755
R404 x9.V2.n121 x9.V2.n112 0.7755
R405 x9.V2.n120 x9.V2.n111 0.7755
R406 x9.V2.n119 x9.V2.n110 0.7755
R407 x9.V2.n118 x9.V2.n109 0.7755
R408 x9.V2.n117 x9.V2.n108 0.7755
R409 x9.V2.n116 x9.V2.n107 0.7755
R410 x9.V2.n106 x9.V2.n2 0.7755
R411 x9.V2.n128 x9.V2.n127 0.7755
R412 x9.V2.n105 x9.V2.n3 0.7755
R413 x9.V2.n104 x9.V2.n103 0.7755
R414 x9.V2.n102 x9.V2.n53 0.7755
R415 x9.V2.n101 x9.V2.n52 0.7755
R416 x9.V2.n100 x9.V2.n51 0.7755
R417 x9.V2.n99 x9.V2.n50 0.7755
R418 x9.V2.n98 x9.V2.n49 0.7755
R419 x9.V2.n97 x9.V2.n48 0.7755
R420 x9.V2.n96 x9.V2.n47 0.7755
R421 x9.V2.n95 x9.V2.n46 0.7755
R422 x9.V2.n94 x9.V2.n45 0.7755
R423 x9.V2.n93 x9.V2.n44 0.7755
R424 x9.V2.n92 x9.V2.n43 0.7755
R425 x9.V2.n91 x9.V2.n42 0.7755
R426 x9.V2.n90 x9.V2.n41 0.7755
R427 x9.V2.n89 x9.V2.n40 0.7755
R428 x9.V2.n88 x9.V2.n39 0.7755
R429 x9.V2.n87 x9.V2.n38 0.7755
R430 x9.V2.n86 x9.V2.n37 0.7755
R431 x9.V2.n85 x9.V2.n36 0.7755
R432 x9.V2.n84 x9.V2.n35 0.7755
R433 x9.V2.n83 x9.V2.n34 0.7755
R434 x9.V2.n82 x9.V2.n33 0.7755
R435 x9.V2.n81 x9.V2.n32 0.7755
R436 x9.V2.n79 x9.V2.n30 0.7755
R437 x9.V2.n78 x9.V2.n29 0.7755
R438 x9.V2.n77 x9.V2.n28 0.7755
R439 x9.V2.n76 x9.V2.n27 0.7755
R440 x9.V2.n75 x9.V2.n26 0.7755
R441 x9.V2.n74 x9.V2.n25 0.7755
R442 x9.V2.n73 x9.V2.n24 0.7755
R443 x9.V2.n72 x9.V2.n23 0.7755
R444 x9.V2.n71 x9.V2.n22 0.7755
R445 x9.V2.n70 x9.V2.n21 0.7755
R446 x9.V2.n69 x9.V2.n20 0.7755
R447 x9.V2.n68 x9.V2.n19 0.7755
R448 x9.V2.n67 x9.V2.n18 0.7755
R449 x9.V2.n66 x9.V2.n17 0.7755
R450 x9.V2.n65 x9.V2.n16 0.7755
R451 x9.V2.n64 x9.V2.n15 0.7755
R452 x9.V2.n63 x9.V2.n14 0.7755
R453 x9.V2.n62 x9.V2.n13 0.7755
R454 x9.V2.n61 x9.V2.n12 0.7755
R455 x9.V2.n60 x9.V2.n11 0.7755
R456 x9.V2.n59 x9.V2.n10 0.7755
R457 x9.V2.n58 x9.V2.n9 0.7755
R458 x9.V2.n57 x9.V2.n8 0.7755
R459 x9.V2.n56 x9.V2.n7 0.7755
R460 x9.V2.n55 x9.V2.n6 0.7755
R461 x9.V2.n54 x9.V2.n5 0.7755
R462 x9.V2.n80 x9.V2.n31 0.7755
R463 x9.V2.n31 x9.V2.t0 0.763824
R464 x9.V2.n126 x9.V2.n4 0.649775
R465 x9.V2.n126 x9.V2.n5 0.649775
R466 x9.V2.n126 x9.V2.n6 0.649775
R467 x9.V2.n126 x9.V2.n7 0.649775
R468 x9.V2.n126 x9.V2.n8 0.649775
R469 x9.V2.n126 x9.V2.n9 0.649775
R470 x9.V2.n126 x9.V2.n10 0.649775
R471 x9.V2.n126 x9.V2.n11 0.649775
R472 x9.V2.n126 x9.V2.n12 0.649775
R473 x9.V2.n126 x9.V2.n13 0.649775
R474 x9.V2.n126 x9.V2.n14 0.649775
R475 x9.V2.n126 x9.V2.n15 0.649775
R476 x9.V2.n126 x9.V2.n16 0.649775
R477 x9.V2.n126 x9.V2.n17 0.649775
R478 x9.V2.n126 x9.V2.n18 0.649775
R479 x9.V2.n126 x9.V2.n19 0.649775
R480 x9.V2.n126 x9.V2.n20 0.649775
R481 x9.V2.n126 x9.V2.n21 0.649775
R482 x9.V2.n126 x9.V2.n22 0.649775
R483 x9.V2.n126 x9.V2.n23 0.649775
R484 x9.V2.n126 x9.V2.n24 0.649775
R485 x9.V2.n126 x9.V2.n25 0.649775
R486 x9.V2.n126 x9.V2.n26 0.649775
R487 x9.V2.n126 x9.V2.n27 0.649775
R488 x9.V2.n126 x9.V2.n28 0.649775
R489 x9.V2.n126 x9.V2.n29 0.649775
R490 x9.V2.n126 x9.V2.n30 0.649775
R491 x9.V2.n126 x9.V2.n31 0.649775
R492 x9.V2.n126 x9.V2.n32 0.649775
R493 x9.V2.n126 x9.V2.n33 0.649775
R494 x9.V2.n126 x9.V2.n34 0.649775
R495 x9.V2.n126 x9.V2.n35 0.649775
R496 x9.V2.n126 x9.V2.n36 0.649775
R497 x9.V2.n126 x9.V2.n37 0.649775
R498 x9.V2.n126 x9.V2.n38 0.649775
R499 x9.V2.n126 x9.V2.n39 0.649775
R500 x9.V2.n126 x9.V2.n40 0.649775
R501 x9.V2.n126 x9.V2.n41 0.649775
R502 x9.V2.n126 x9.V2.n42 0.649775
R503 x9.V2.n126 x9.V2.n43 0.649775
R504 x9.V2.n126 x9.V2.n44 0.649775
R505 x9.V2.n126 x9.V2.n45 0.649775
R506 x9.V2.n126 x9.V2.n46 0.649775
R507 x9.V2.n126 x9.V2.n47 0.649775
R508 x9.V2.n126 x9.V2.n48 0.649775
R509 x9.V2.n126 x9.V2.n49 0.649775
R510 x9.V2.n126 x9.V2.n50 0.649775
R511 x9.V2.n126 x9.V2.n51 0.649775
R512 x9.V2.n126 x9.V2.n52 0.649775
R513 x9.V2.n126 x9.V2.n53 0.649775
R514 x9.V2.n126 x9.V2.n104 0.649775
R515 x9.V2.n126 x9.V2.n105 0.649775
R516 x9.V2.n127 x9.V2.n126 0.649775
R517 x9.V2.n126 x9.V2.n106 0.649775
R518 x9.V2.n126 x9.V2.n107 0.649775
R519 x9.V2.n126 x9.V2.n108 0.649775
R520 x9.V2.n126 x9.V2.n109 0.649775
R521 x9.V2.n126 x9.V2.n110 0.649775
R522 x9.V2.n126 x9.V2.n111 0.649775
R523 x9.V2.n126 x9.V2.n112 0.649775
R524 x9.V2.n126 x9.V2.n113 0.649775
R525 x9.V2.n126 x9.V2.n114 0.649775
R526 x9.V2.n126 x9.V2.n115 0.649775
R527 x9.V2.n126 x9.V2.n125 0.649775
R528 x9.V2 x9.V2.n137 0.399458
R529 x9.V2.n134 x9.V2.n133 0.219746
R530 x9.V2.n136 x9.V2.n134 0.0892897
R531 x9.V2.n124 x9.V2.n123 0.068052
R532 x9.V2.n123 x9.V2.n122 0.068052
R533 x9.V2.n122 x9.V2.n121 0.068052
R534 x9.V2.n121 x9.V2.n120 0.068052
R535 x9.V2.n120 x9.V2.n119 0.068052
R536 x9.V2.n119 x9.V2.n118 0.068052
R537 x9.V2.n118 x9.V2.n117 0.068052
R538 x9.V2.n117 x9.V2.n116 0.068052
R539 x9.V2.n116 x9.V2.n2 0.068052
R540 x9.V2.n128 x9.V2.n3 0.068052
R541 x9.V2.n103 x9.V2.n3 0.068052
R542 x9.V2.n103 x9.V2.n102 0.068052
R543 x9.V2.n102 x9.V2.n101 0.068052
R544 x9.V2.n101 x9.V2.n100 0.068052
R545 x9.V2.n100 x9.V2.n99 0.068052
R546 x9.V2.n99 x9.V2.n98 0.068052
R547 x9.V2.n98 x9.V2.n97 0.068052
R548 x9.V2.n97 x9.V2.n96 0.068052
R549 x9.V2.n96 x9.V2.n95 0.068052
R550 x9.V2.n95 x9.V2.n94 0.068052
R551 x9.V2.n94 x9.V2.n93 0.068052
R552 x9.V2.n93 x9.V2.n92 0.068052
R553 x9.V2.n92 x9.V2.n91 0.068052
R554 x9.V2.n91 x9.V2.n90 0.068052
R555 x9.V2.n90 x9.V2.n89 0.068052
R556 x9.V2.n89 x9.V2.n88 0.068052
R557 x9.V2.n88 x9.V2.n87 0.068052
R558 x9.V2.n87 x9.V2.n86 0.068052
R559 x9.V2.n86 x9.V2.n85 0.068052
R560 x9.V2.n85 x9.V2.n84 0.068052
R561 x9.V2.n84 x9.V2.n83 0.068052
R562 x9.V2.n83 x9.V2.n82 0.068052
R563 x9.V2.n82 x9.V2.n81 0.068052
R564 x9.V2.n81 x9.V2.n80 0.068052
R565 x9.V2.n80 x9.V2.n79 0.068052
R566 x9.V2.n79 x9.V2.n78 0.068052
R567 x9.V2.n78 x9.V2.n77 0.068052
R568 x9.V2.n77 x9.V2.n76 0.068052
R569 x9.V2.n76 x9.V2.n75 0.068052
R570 x9.V2.n75 x9.V2.n74 0.068052
R571 x9.V2.n74 x9.V2.n73 0.068052
R572 x9.V2.n73 x9.V2.n72 0.068052
R573 x9.V2.n72 x9.V2.n71 0.068052
R574 x9.V2.n71 x9.V2.n70 0.068052
R575 x9.V2.n70 x9.V2.n69 0.068052
R576 x9.V2.n69 x9.V2.n68 0.068052
R577 x9.V2.n68 x9.V2.n67 0.068052
R578 x9.V2.n67 x9.V2.n66 0.068052
R579 x9.V2.n66 x9.V2.n65 0.068052
R580 x9.V2.n65 x9.V2.n64 0.068052
R581 x9.V2.n64 x9.V2.n63 0.068052
R582 x9.V2.n63 x9.V2.n62 0.068052
R583 x9.V2.n62 x9.V2.n61 0.068052
R584 x9.V2.n61 x9.V2.n60 0.068052
R585 x9.V2.n60 x9.V2.n59 0.068052
R586 x9.V2.n59 x9.V2.n58 0.068052
R587 x9.V2.n58 x9.V2.n57 0.068052
R588 x9.V2.n57 x9.V2.n56 0.068052
R589 x9.V2.n56 x9.V2.n55 0.068052
R590 x9.V2.n55 x9.V2.n54 0.068052
R591 x9.V2.n129 x9.V2.n128 0.0417818
R592 x9.V2.n129 x9.V2.n2 0.0267702
R593 VSS.n893 VSS.n892 6.38338e+06
R594 VSS.n1252 VSS.n244 134296
R595 VSS.n916 VSS.n540 53810
R596 VSS.n896 VSS.n540 53810
R597 VSS.n894 VSS.n557 53810
R598 VSS.n914 VSS.n557 53810
R599 VSS.n904 VSS.n575 43763
R600 VSS.n904 VSS.n539 43763
R601 VSS.n906 VSS.n574 43763
R602 VSS.n906 VSS.n558 43763
R603 VSS.n1104 VSS.n408 21270.2
R604 VSS.n1089 VSS.n408 21270.2
R605 VSS.n1104 VSS.n409 21270.2
R606 VSS.n1089 VSS.n409 21270.2
R607 VSS.n944 VSS.n534 21270.2
R608 VSS.n944 VSS.n11 21270.2
R609 VSS.n534 VSS.n532 21270.2
R610 VSS.n532 VSS.n11 21270.2
R611 VSS.n1106 VSS.n407 21270.2
R612 VSS.n407 VSS.n394 21270.2
R613 VSS.n1107 VSS.n1106 21270.2
R614 VSS.n1107 VSS.n394 21270.2
R615 VSS.n533 VSS.n529 21270.2
R616 VSS.n533 VSS.n530 21270.2
R617 VSS.n946 VSS.n529 21270.2
R618 VSS.n946 VSS.n530 21270.2
R619 VSS.n374 VSS.n373 15846.9
R620 VSS.n1132 VSS.n373 15846.9
R621 VSS.n1131 VSS.n374 15846.9
R622 VSS.n1132 VSS.n1131 15846.9
R623 VSS.n1436 VSS.n8 15846.9
R624 VSS.n1418 VSS.n8 15846.9
R625 VSS.n1436 VSS.n9 15846.9
R626 VSS.n1418 VSS.n9 15846.9
R627 VSS.n369 VSS.n368 15846.9
R628 VSS.n1134 VSS.n369 15846.9
R629 VSS.n1135 VSS.n368 15846.9
R630 VSS.n1135 VSS.n1134 15846.9
R631 VSS.n34 VSS.n6 15846.9
R632 VSS.n1420 VSS.n34 15846.9
R633 VSS.n1421 VSS.n6 15846.9
R634 VSS.n1421 VSS.n1420 15846.9
R635 VSS.n182 VSS.n181 13135.3
R636 VSS.n1303 VSS.n182 13135.3
R637 VSS.n1304 VSS.n181 13135.3
R638 VSS.n1304 VSS.n1303 13135.3
R639 VSS.n728 VSS.n58 13135.3
R640 VSS.n1401 VSS.n58 13135.3
R641 VSS.n728 VSS.n59 13135.3
R642 VSS.n1401 VSS.n59 13135.3
R643 VSS.n762 VSS.n742 13135.3
R644 VSS.n742 VSS.n185 13135.3
R645 VSS.n762 VSS.n743 13135.3
R646 VSS.n743 VSS.n185 13135.3
R647 VSS.n56 VSS.n55 13135.3
R648 VSS.n1403 VSS.n56 13135.3
R649 VSS.n1404 VSS.n55 13135.3
R650 VSS.n1404 VSS.n1403 13135.3
R651 VSS.n327 VSS.n280 11779.4
R652 VSS.n1212 VSS.n280 11779.4
R653 VSS.n327 VSS.n281 11779.4
R654 VSS.n1212 VSS.n281 11779.4
R655 VSS.n792 VSS.n81 11779.4
R656 VSS.n1384 VSS.n81 11779.4
R657 VSS.n792 VSS.n82 11779.4
R658 VSS.n1384 VSS.n82 11779.4
R659 VSS.n277 VSS.n276 11779.4
R660 VSS.n1214 VSS.n277 11779.4
R661 VSS.n1215 VSS.n276 11779.4
R662 VSS.n1215 VSS.n1214 11779.4
R663 VSS.n78 VSS.n77 11779.4
R664 VSS.n1386 VSS.n78 11779.4
R665 VSS.n1387 VSS.n77 11779.4
R666 VSS.n1387 VSS.n1386 11779.4
R667 VSS.n311 VSS.n221 11101.5
R668 VSS.n1272 VSS.n221 11101.5
R669 VSS.n311 VSS.n222 11101.5
R670 VSS.n1272 VSS.n222 11101.5
R671 VSS.n1210 VSS.n283 11101.5
R672 VSS.n313 VSS.n283 11101.5
R673 VSS.n1210 VSS.n314 11101.5
R674 VSS.n314 VSS.n313 11101.5
R675 VSS.n1039 VSS.n461 11101.5
R676 VSS.n1039 VSS.n462 11101.5
R677 VSS.n461 VSS.n460 11101.5
R678 VSS.n462 VSS.n460 11101.5
R679 VSS.n1382 VSS.n84 11101.5
R680 VSS.n483 VSS.n84 11101.5
R681 VSS.n1382 VSS.n85 11101.5
R682 VSS.n483 VSS.n85 11101.5
R683 VSS.n1180 VSS.n218 11101.5
R684 VSS.n1274 VSS.n218 11101.5
R685 VSS.n1180 VSS.n219 11101.5
R686 VSS.n1274 VSS.n219 11101.5
R687 VSS.n1172 VSS.n316 11101.5
R688 VSS.n1182 VSS.n1172 11101.5
R689 VSS.n1183 VSS.n316 11101.5
R690 VSS.n1183 VSS.n1182 11101.5
R691 VSS.n458 VSS.n457 11101.5
R692 VSS.n1041 VSS.n457 11101.5
R693 VSS.n1040 VSS.n458 11101.5
R694 VSS.n1041 VSS.n1040 11101.5
R695 VSS.n1002 VSS.n87 11101.5
R696 VSS.n1005 VSS.n1002 11101.5
R697 VSS.n1004 VSS.n87 11101.5
R698 VSS.n1005 VSS.n1004 11101.5
R699 VSS.n916 VSS.n539 10047
R700 VSS.n591 VSS.n574 10047
R701 VSS.n591 VSS.n575 10047
R702 VSS.n896 VSS.n575 10047
R703 VSS.n894 VSS.n574 10047
R704 VSS.n914 VSS.n558 10047
R705 VSS.n558 VSS.n541 10047
R706 VSS.n541 VSS.n539 10047
R707 VSS.n1094 VSS.n426 8377.66
R708 VSS.n436 VSS.n426 8377.66
R709 VSS.n436 VSS.n422 8377.66
R710 VSS.n1094 VSS.n422 8377.66
R711 VSS.n626 VSS.n621 8377.66
R712 VSS.n627 VSS.n621 8377.66
R713 VSS.n666 VSS.n627 8377.66
R714 VSS.n666 VSS.n626 8377.66
R715 VSS.n1092 VSS.n1091 8377.66
R716 VSS.n1091 VSS.n437 8377.66
R717 VSS.n1059 VSS.n437 8377.66
R718 VSS.n1092 VSS.n1059 8377.66
R719 VSS.n691 VSS.n622 8377.66
R720 VSS.n691 VSS.n623 8377.66
R721 VSS.n668 VSS.n623 8377.66
R722 VSS.n668 VSS.n622 8377.66
R723 VSS.n551 VSS.n542 7765.14
R724 VSS.n551 VSS.n544 7765.14
R725 VSS.n555 VSS.n544 7765.14
R726 VSS.n555 VSS.n542 7765.14
R727 VSS.n891 VSS.n594 7663.05
R728 VSS.n594 VSS.n592 7663.05
R729 VSS.n593 VSS.n592 7663.05
R730 VSS.n891 VSS.n593 7663.05
R731 VSS.n249 VSS.n171 7663.05
R732 VSS.n249 VSS.n172 7663.05
R733 VSS.n1310 VSS.n172 7663.05
R734 VSS.n1310 VSS.n171 7663.05
R735 VSS.n1064 VSS.n130 7663.05
R736 VSS.n1064 VSS.n131 7663.05
R737 VSS.n1343 VSS.n131 7663.05
R738 VSS.n1343 VSS.n130 7663.05
R739 VSS.n1362 VSS.n106 7663.05
R740 VSS.n1362 VSS.n107 7663.05
R741 VSS.n1365 VSS.n107 7663.05
R742 VSS.n1365 VSS.n106 7663.05
R743 VSS.n795 VSS.n733 7663.05
R744 VSS.n795 VSS.n734 7663.05
R745 VSS.n827 VSS.n734 7663.05
R746 VSS.n827 VSS.n733 7663.05
R747 VSS.n860 VSS.n695 7663.05
R748 VSS.n696 VSS.n695 7663.05
R749 VSS.n860 VSS.n859 7663.05
R750 VSS.n859 VSS.n696 7663.05
R751 VSS.n873 VSS.n613 6737.69
R752 VSS.n873 VSS.n612 6737.69
R753 VSS.n865 VSS.n620 6737.69
R754 VSS.n866 VSS.n620 6737.69
R755 VSS.n342 VSS.n321 6737.69
R756 VSS.n321 VSS.n320 6737.69
R757 VSS.n1255 VSS.n1254 6737.69
R758 VSS.n1254 VSS.n241 6737.69
R759 VSS.n1321 VSS.n161 6737.69
R760 VSS.n1320 VSS.n161 6737.69
R761 VSS.n1316 VSS.n167 6737.69
R762 VSS.n1315 VSS.n167 6737.69
R763 VSS.n1349 VSS.n123 6737.69
R764 VSS.n1349 VSS.n124 6737.69
R765 VSS.n1339 VSS.n136 6737.69
R766 VSS.n1338 VSS.n136 6737.69
R767 VSS.n1376 VSS.n94 6737.69
R768 VSS.n1375 VSS.n94 6737.69
R769 VSS.n1371 VSS.n101 6737.69
R770 VSS.n1370 VSS.n101 6737.69
R771 VSS.n838 VSS.n720 6737.69
R772 VSS.n837 VSS.n720 6737.69
R773 VSS.n833 VSS.n727 6737.69
R774 VSS.n832 VSS.n727 6737.69
R775 VSS.n878 VSS.n605 6490.71
R776 VSS.n887 VSS.n598 6490.71
R777 VSS.n887 VSS.n884 6490.71
R778 VSS.n879 VSS.n605 6490.71
R779 VSS.n1300 VSS.n189 6490.71
R780 VSS.n189 VSS.n188 6490.71
R781 VSS.n338 VSS.n337 6490.71
R782 VSS.n338 VSS.n323 6490.71
R783 VSS.n1332 VSS.n145 6490.71
R784 VSS.n1331 VSS.n145 6490.71
R785 VSS.n1326 VSS.n152 6490.71
R786 VSS.n1325 VSS.n152 6490.71
R787 VSS.n432 VSS.n431 6490.71
R788 VSS.n431 VSS.n429 6490.71
R789 VSS.n1353 VSS.n117 6490.71
R790 VSS.n1354 VSS.n117 6490.71
R791 VSS.n800 VSS.n788 6490.71
R792 VSS.n801 VSS.n788 6490.71
R793 VSS.n90 VSS.n88 6490.71
R794 VSS.n1380 VSS.n90 6490.71
R795 VSS.n842 VSS.n713 6490.71
R796 VSS.n856 VSS.n697 6490.71
R797 VSS.n856 VSS.n698 6490.71
R798 VSS.n843 VSS.n713 6490.71
R799 VSS.n332 VSS.n245 5875.23
R800 VSS.n1251 VSS.n245 5875.23
R801 VSS.n332 VSS.n246 5875.23
R802 VSS.n1251 VSS.n246 5875.23
R803 VSS.n769 VSS.n150 5875.23
R804 VSS.n769 VSS.n766 5875.23
R805 VSS.n770 VSS.n150 5875.23
R806 VSS.n770 VSS.n766 5875.23
R807 VSS.n1347 VSS.n127 5875.23
R808 VSS.n1347 VSS.n1346 5875.23
R809 VSS.n127 VSS.n126 5875.23
R810 VSS.n1346 VSS.n126 5875.23
R811 VSS.n809 VSS.n808 5875.23
R812 VSS.n813 VSS.n809 5875.23
R813 VSS.n814 VSS.n808 5875.23
R814 VSS.n814 VSS.n813 5875.23
R815 VSS.n846 VSS.n710 5875.23
R816 VSS.n824 VSS.n710 5875.23
R817 VSS.n846 VSS.n711 5875.23
R818 VSS.n824 VSS.n711 5875.23
R819 VSS.n603 VSS.n3 5875.23
R820 VSS.n603 VSS.n4 5875.23
R821 VSS.n1439 VSS.n3 5875.23
R822 VSS.n1439 VSS.n4 5875.23
R823 VSS.n1126 VSS.n378 5822.21
R824 VSS.n1126 VSS.n1125 5822.21
R825 VSS.n1125 VSS.n379 5822.21
R826 VSS.n379 VSS.n378 5822.21
R827 VSS.n1426 VSS.n26 5822.21
R828 VSS.n27 VSS.n26 5822.21
R829 VSS.n27 VSS.n25 5822.21
R830 VSS.n1426 VSS.n25 5822.21
R831 VSS.n1139 VSS.n1138 5822.21
R832 VSS.n1140 VSS.n1139 5822.21
R833 VSS.n1140 VSS.n363 5822.21
R834 VSS.n1138 VSS.n363 5822.21
R835 VSS.n1424 VSS.n31 5822.21
R836 VSS.n31 VSS.n28 5822.21
R837 VSS.n30 VSS.n28 5822.21
R838 VSS.n1424 VSS.n30 5822.21
R839 VSS.n870 VSS.n615 5089.59
R840 VSS.n870 VSS.n616 5089.59
R841 VSS.n1259 VSS.n236 5089.59
R842 VSS.n1259 VSS.n237 5089.59
R843 VSS.n371 VSS.n162 5089.59
R844 VSS.n371 VSS.n163 5089.59
R845 VSS.n139 VSS.n137 5089.59
R846 VSS.n139 VSS.n135 5089.59
R847 VSS.n102 VSS.n95 5089.59
R848 VSS.n102 VSS.n97 5089.59
R849 VSS.n730 VSS.n721 5089.59
R850 VSS.n730 VSS.n723 5089.59
R851 VSS.n609 VSS.n608 4951.75
R852 VSS.n329 VSS.n190 4951.75
R853 VSS.n153 VSS.n146 4951.75
R854 VSS.n433 VSS.n116 4951.75
R855 VSS.n805 VSS.n89 4951.75
R856 VSS.n849 VSS.n708 4951.75
R857 VSS.n608 VSS.n599 4948.9
R858 VSS.n329 VSS.n324 4948.9
R859 VSS.n153 VSS.n147 4948.9
R860 VSS.n433 VSS.n119 4948.9
R861 VSS.n805 VSS.n785 4948.9
R862 VSS.n849 VSS.n709 4948.9
R863 VSS.n1307 VSS.n178 4211.88
R864 VSS.n178 VSS.n173 4211.88
R865 VSS.n177 VSS.n173 4211.88
R866 VSS.n1307 VSS.n177 4211.88
R867 VSS.n1409 VSS.n47 4211.88
R868 VSS.n48 VSS.n47 4211.88
R869 VSS.n48 VSS.n46 4211.88
R870 VSS.n1409 VSS.n46 4211.88
R871 VSS.n186 VSS.n176 4211.88
R872 VSS.n186 VSS.n174 4211.88
R873 VSS.n365 VSS.n174 4211.88
R874 VSS.n365 VSS.n176 4211.88
R875 VSS.n1407 VSS.n52 4211.88
R876 VSS.n52 VSS.n49 4211.88
R877 VSS.n51 VSS.n49 4211.88
R878 VSS.n1407 VSS.n51 4211.88
R879 VSS.n1220 VSS.n268 3434.71
R880 VSS.n269 VSS.n268 3434.71
R881 VSS.n269 VSS.n267 3434.71
R882 VSS.n1220 VSS.n267 3434.71
R883 VSS.n1392 VSS.n69 3434.71
R884 VSS.n70 VSS.n69 3434.71
R885 VSS.n70 VSS.n68 3434.71
R886 VSS.n1392 VSS.n68 3434.71
R887 VSS.n1218 VSS.n273 3434.71
R888 VSS.n273 VSS.n270 3434.71
R889 VSS.n272 VSS.n270 3434.71
R890 VSS.n1218 VSS.n272 3434.71
R891 VSS.n1390 VSS.n74 3434.71
R892 VSS.n74 VSS.n71 3434.71
R893 VSS.n73 VSS.n71 3434.71
R894 VSS.n1390 VSS.n73 3434.71
R895 VSS.n1050 VSS.n411 3175.68
R896 VSS.n210 VSS.n200 3153.92
R897 VSS.n1208 VSS.n344 2976.97
R898 VSS.n344 VSS.n343 2976.97
R899 VSS.n207 VSS.n205 2976.97
R900 VSS.n1288 VSS.n207 2976.97
R901 VSS.n998 VSS.n993 2976.97
R902 VSS.n999 VSS.n998 2976.97
R903 VSS.n1051 VSS.n445 2976.97
R904 VSS.n1051 VSS.n444 2976.97
R905 VSS.n1147 VSS.n318 2976.97
R906 VSS.n1147 VSS.n319 2976.97
R907 VSS.n1289 VSS.n203 2976.97
R908 VSS.n204 VSS.n203 2976.97
R909 VSS.n679 VSS.n678 2976.97
R910 VSS.n680 VSS.n679 2976.97
R911 VSS.n1054 VSS.n1053 2976.97
R912 VSS.n1053 VSS.n443 2976.97
R913 VSS.n1283 VSS.n210 2410.42
R914 VSS.n1292 VSS.n1291 2011.1
R915 VSS.n1262 VSS.n206 1881.91
R916 VSS.n1262 VSS.n232 1881.91
R917 VSS.n1018 VSS.n493 1881.91
R918 VSS.n1018 VSS.n494 1881.91
R919 VSS.n317 VSS.n234 1881.91
R920 VSS.n234 VSS.n202 1881.91
R921 VSS.n1014 VSS.n496 1881.91
R922 VSS.n1014 VSS.n442 1881.91
R923 VSS.n908 VSS.n907 1663.12
R924 VSS.n907 VSS.n573 1663.12
R925 VSS.n1292 VSS.n199 1151.27
R926 VSS.n920 VSS.n535 1061.93
R927 VSS.n922 VSS.n535 1004.8
R928 VSS.n566 VSS.n561 975.168
R929 VSS.n568 VSS.n567 975.168
R930 VSS.n569 VSS.n559 975.168
R931 VSS.n912 VSS.n911 975.168
R932 VSS.n910 VSS.n560 975.168
R933 VSS.n909 VSS.n571 975.168
R934 VSS.n584 VSS.n582 975.105
R935 VSS.n585 VSS.n579 975.105
R936 VSS.n589 VSS.n588 975.105
R937 VSS.n587 VSS.n581 975.105
R938 VSS.n580 VSS.n577 975.105
R939 VSS.n583 VSS.n572 975.105
R940 VSS.n919 VSS.n536 969.856
R941 VSS.n918 VSS.n537 969.856
R942 VSS.n898 VSS.n538 969.856
R943 VSS.n900 VSS.n899 969.856
R944 VSS.n901 VSS.n578 969.856
R945 VSS.n921 VSS.n920 969.856
R946 VSS.n923 VSS.n922 946.241
R947 VSS.n903 VSS.n576 910.009
R948 VSS.n903 VSS.n902 910.009
R949 VSS.n890 VSS.n595 819.808
R950 VSS.n600 VSS.n595 816.99
R951 VSS.n884 VSS.n599 773.438
R952 VSS.n324 VSS.n188 773.438
R953 VSS.n1331 VSS.n147 773.438
R954 VSS.n429 VSS.n119 773.438
R955 VSS.n801 VSS.n785 773.438
R956 VSS.n709 VSS.n698 773.438
R957 VSS.n878 VSS.n609 770.587
R958 VSS.n609 VSS.n598 770.587
R959 VSS.n879 VSS.n599 770.587
R960 VSS.n616 VSS.n613 770.587
R961 VSS.n865 VSS.n615 770.587
R962 VSS.n615 VSS.n612 770.587
R963 VSS.n866 VSS.n616 770.587
R964 VSS.n1300 VSS.n190 770.587
R965 VSS.n337 VSS.n324 770.587
R966 VSS.n323 VSS.n190 770.587
R967 VSS.n342 VSS.n236 770.587
R968 VSS.n320 VSS.n237 770.587
R969 VSS.n1255 VSS.n237 770.587
R970 VSS.n241 VSS.n236 770.587
R971 VSS.n1332 VSS.n146 770.587
R972 VSS.n1326 VSS.n147 770.587
R973 VSS.n1325 VSS.n146 770.587
R974 VSS.n1321 VSS.n162 770.587
R975 VSS.n1320 VSS.n163 770.587
R976 VSS.n1316 VSS.n163 770.587
R977 VSS.n1315 VSS.n162 770.587
R978 VSS.n432 VSS.n116 770.587
R979 VSS.n1353 VSS.n119 770.587
R980 VSS.n1354 VSS.n116 770.587
R981 VSS.n137 VSS.n123 770.587
R982 VSS.n135 VSS.n124 770.587
R983 VSS.n1339 VSS.n135 770.587
R984 VSS.n1338 VSS.n137 770.587
R985 VSS.n800 VSS.n89 770.587
R986 VSS.n785 VSS.n88 770.587
R987 VSS.n1380 VSS.n89 770.587
R988 VSS.n1376 VSS.n95 770.587
R989 VSS.n1375 VSS.n97 770.587
R990 VSS.n1371 VSS.n97 770.587
R991 VSS.n1370 VSS.n95 770.587
R992 VSS.n842 VSS.n708 770.587
R993 VSS.n708 VSS.n697 770.587
R994 VSS.n843 VSS.n709 770.587
R995 VSS.n838 VSS.n721 770.587
R996 VSS.n837 VSS.n723 770.587
R997 VSS.n833 VSS.n723 770.587
R998 VSS.n832 VSS.n721 770.587
R999 VSS.n1208 VSS.n206 770.587
R1000 VSS.n343 VSS.n232 770.587
R1001 VSS.n232 VSS.n205 770.587
R1002 VSS.n1288 VSS.n206 770.587
R1003 VSS.n993 VSS.n493 770.587
R1004 VSS.n999 VSS.n494 770.587
R1005 VSS.n494 VSS.n445 770.587
R1006 VSS.n493 VSS.n444 770.587
R1007 VSS.n318 VSS.n317 770.587
R1008 VSS.n319 VSS.n202 770.587
R1009 VSS.n1289 VSS.n202 770.587
R1010 VSS.n317 VSS.n204 770.587
R1011 VSS.n678 VSS.n496 770.587
R1012 VSS.n680 VSS.n442 770.587
R1013 VSS.n1054 VSS.n442 770.587
R1014 VSS.n496 VSS.n443 770.587
R1015 VSS.n1080 VSS.n1078 652.918
R1016 VSS.n1318 VSS.n165 522.183
R1017 VSS.n140 VSS.n134 522.183
R1018 VSS.n1373 VSS.n99 522.183
R1019 VSS.n835 VSS.n725 522.183
R1020 VSS.n1258 VSS.n1257 522.183
R1021 VSS.n869 VSS.n868 522.183
R1022 VSS.n165 VSS.n159 509.091
R1023 VSS.n142 VSS.n140 509.091
R1024 VSS.n99 VSS.n93 509.091
R1025 VSS.n725 VSS.n718 509.091
R1026 VSS.n1258 VSS.n238 509.091
R1027 VSS.n869 VSS.n617 509.091
R1028 VSS.n1110 VSS.n405 494.08
R1029 VSS.n1111 VSS.n403 494.08
R1030 VSS.n1112 VSS.n401 494.08
R1031 VSS.n1113 VSS.n399 494.08
R1032 VSS.n1114 VSS.n397 494.08
R1033 VSS.n1117 VSS.n391 494.08
R1034 VSS.n1118 VSS.n389 494.08
R1035 VSS.n1119 VSS.n387 494.08
R1036 VSS.n1120 VSS.n385 494.08
R1037 VSS.n1121 VSS.n383 494.08
R1038 VSS.n1116 VSS.n393 493.697
R1039 VSS.n1097 VSS.n419 491.521
R1040 VSS.n1098 VSS.n418 491.521
R1041 VSS.n1099 VSS.n414 491.521
R1042 VSS.n1100 VSS.n413 491.521
R1043 VSS.n1101 VSS.n412 491.521
R1044 VSS.n1087 VSS.n410 491.521
R1045 VSS.n1086 VSS.n1070 491.521
R1046 VSS.n1085 VSS.n1072 491.521
R1047 VSS.n1084 VSS.n1074 491.521
R1048 VSS.n1083 VSS.n1076 491.521
R1049 VSS.n1082 VSS.n1078 491.521
R1050 VSS.n949 VSS.n527 491.521
R1051 VSS.n653 VSS.n526 491.521
R1052 VSS.n654 VSS.n525 491.521
R1053 VSS.n655 VSS.n524 491.521
R1054 VSS.n656 VSS.n523 491.521
R1055 VSS.n658 VSS.n652 491.521
R1056 VSS.n659 VSS.n635 491.521
R1057 VSS.n660 VSS.n634 491.521
R1058 VSS.n661 VSS.n633 491.521
R1059 VSS.n662 VSS.n632 491.521
R1060 VSS.n663 VSS.n631 491.521
R1061 VSS.n1430 VSS.n21 491.521
R1062 VSS.n1431 VSS.n19 491.521
R1063 VSS.n1432 VSS.n17 491.521
R1064 VSS.n1433 VSS.n15 491.521
R1065 VSS.n1434 VSS.n13 491.521
R1066 VSS.n935 VSS.n10 491.521
R1067 VSS.n937 VSS.n936 491.521
R1068 VSS.n938 VSS.n932 491.521
R1069 VSS.n939 VSS.n930 491.521
R1070 VSS.n940 VSS.n928 491.521
R1071 VSS.n941 VSS.n926 491.521
R1072 VSS.n563 VSS.n562 456.122
R1073 VSS.n1081 VSS.n1080 431.159
R1074 VSS.n243 VSS.n242 418.079
R1075 VSS.n243 VSS.n240 410.286
R1076 VSS.n553 VSS.n552 382.872
R1077 VSS.n554 VSS.n553 380.592
R1078 VSS.n1050 VSS 348.952
R1079 VSS.n1250 VSS.n1249 338.159
R1080 VSS.n1057 VSS.n1055 312.123
R1081 VSS.n1248 VSS.n251 305.545
R1082 VSS.n565 VSS.n564 303.812
R1083 VSS.n564 VSS.n563 303.772
R1084 VSS.n499 VSS.n440 298.668
R1085 VSS.n772 VSS.n148 295.589
R1086 VSS.n777 VSS.n109 295.589
R1087 VSS.n816 VSS.n737 295.589
R1088 VSS.n820 VSS.n700 295.589
R1089 VSS.n915 VSS.n556 294.541
R1090 VSS.n815 VSS.n780 290.49
R1091 VSS.n776 VSS.n775 290.49
R1092 VSS.n771 VSS.n740 290.49
R1093 VSS.n822 VSS.n821 290.49
R1094 VSS.n1097 VSS.n1096 286.08
R1095 VSS.n1329 VSS.n149 280.81
R1096 VSS.n427 VSS.n112 280.81
R1097 VSS.n804 VSS.n803 280.81
R1098 VSS.n326 VSS.n193 280.81
R1099 VSS.n850 VSS.n707 280.81
R1100 VSS.n882 VSS.n602 280.81
R1101 VSS.n1096 VSS.n420 268.387
R1102 VSS.n562 VSS.n199 265.623
R1103 VSS.n1110 VSS.n404 251.905
R1104 VSS.n1111 VSS.n402 251.905
R1105 VSS.n1112 VSS.n400 251.905
R1106 VSS.n1113 VSS.n398 251.905
R1107 VSS.n1114 VSS.n395 251.905
R1108 VSS.n1116 VSS.n392 251.905
R1109 VSS.n1117 VSS.n390 251.905
R1110 VSS.n1118 VSS.n388 251.905
R1111 VSS.n1119 VSS.n386 251.905
R1112 VSS.n1120 VSS.n384 251.905
R1113 VSS.n1121 VSS.n382 251.905
R1114 VSS.n419 VSS.n376 251.905
R1115 VSS.n418 VSS.n417 251.905
R1116 VSS.n416 VSS.n414 251.905
R1117 VSS.n415 VSS.n413 251.905
R1118 VSS.n412 VSS.n261 251.905
R1119 VSS.n1087 VSS.n1068 251.905
R1120 VSS.n1086 VSS.n1069 251.905
R1121 VSS.n1085 VSS.n1071 251.905
R1122 VSS.n1084 VSS.n1073 251.905
R1123 VSS.n1083 VSS.n1075 251.905
R1124 VSS.n1082 VSS.n1077 251.905
R1125 VSS.n1430 VSS.n20 251.905
R1126 VSS.n1431 VSS.n18 251.905
R1127 VSS.n1432 VSS.n16 251.905
R1128 VSS.n1433 VSS.n14 251.905
R1129 VSS.n1434 VSS.n12 251.905
R1130 VSS.n38 VSS.n10 251.905
R1131 VSS.n937 VSS.n933 251.905
R1132 VSS.n938 VSS.n931 251.905
R1133 VSS.n939 VSS.n929 251.905
R1134 VSS.n940 VSS.n927 251.905
R1135 VSS.n941 VSS.n925 251.905
R1136 VSS.n950 VSS.n949 251.905
R1137 VSS.n951 VSS.n526 251.905
R1138 VSS.n952 VSS.n525 251.905
R1139 VSS.n953 VSS.n524 251.905
R1140 VSS.n954 VSS.n523 251.905
R1141 VSS.n652 VSS.n650 251.905
R1142 VSS.n649 VSS.n635 251.905
R1143 VSS.n648 VSS.n634 251.905
R1144 VSS.n647 VSS.n633 251.905
R1145 VSS.n646 VSS.n632 251.905
R1146 VSS.n645 VSS.n631 251.905
R1147 VSS.n1050 VSS.n1049 251.798
R1148 VSS.n1079 VSS.n1077 251.346
R1149 VSS.n925 VSS.n924 251.346
R1150 VSS.n438 VSS.n405 233.601
R1151 VSS.n446 VSS.n420 232.18
R1152 VSS.n1081 VSS.n1079 220.969
R1153 VSS.n942 VSS.n924 220.969
R1154 VSS.n446 VSS.n383 204.161
R1155 VSS.n1248 VSS.n1247 200.084
R1156 VSS.n817 VSS.n816 196.312
R1157 VSS.n778 VSS.n777 196.312
R1158 VSS.n773 VSS.n772 196.312
R1159 VSS.n820 VSS.n0 196.312
R1160 VSS.n1328 VSS.n150 195.001
R1161 VSS.n127 VSS.n120 195.001
R1162 VSS.n808 VSS.n784 195.001
R1163 VSS.n333 VSS.n332 195.001
R1164 VSS.n846 VSS.n845 195.001
R1165 VSS.n881 VSS.n603 195.001
R1166 VSS.n1004 VSS.n497 195
R1167 VSS.n1004 VSS.t149 195
R1168 VSS.n1002 VSS.n1001 195
R1169 VSS.t149 VSS.n1002 195
R1170 VSS.n1040 VSS.n459 195
R1171 VSS.n1040 VSS.t106 195
R1172 VSS.n491 VSS.n457 195
R1173 VSS.t106 VSS.n457 195
R1174 VSS.n1184 VSS.n1183 195
R1175 VSS.n1183 VSS.t122 195
R1176 VSS.n1172 VSS.n1171 195
R1177 VSS.n1172 VSS.t122 195
R1178 VSS.n1169 VSS.n219 195
R1179 VSS.n219 VSS.t163 195
R1180 VSS.n230 VSS.n218 195
R1181 VSS.n218 VSS.t163 195
R1182 VSS.n489 VSS.n85 195
R1183 VSS.t149 VSS.n85 195
R1184 VSS.n474 VSS.n84 195
R1185 VSS.t149 VSS.n84 195
R1186 VSS.n1022 VSS.n460 195
R1187 VSS.t106 VSS.n460 195
R1188 VSS.n1039 VSS.n1038 195
R1189 VSS.t106 VSS.n1039 195
R1190 VSS.n314 VSS.n229 195
R1191 VSS.t122 VSS.n314 195
R1192 VSS.n303 VSS.n283 195
R1193 VSS.t122 VSS.n283 195
R1194 VSS.n222 VSS.n208 195
R1195 VSS.n222 VSS.t163 195
R1196 VSS.n294 VSS.n221 195
R1197 VSS.n221 VSS.t163 195
R1198 VSS.n824 VSS.n823 195
R1199 VSS.n825 VSS.n824 195
R1200 VSS.n813 VSS.n810 195
R1201 VSS.n813 VSS.n812 195
R1202 VSS.n808 VSS.n807 195
R1203 VSS.n1346 VSS.n128 195
R1204 VSS.n1346 VSS.n1345 195
R1205 VSS.n435 VSS.n127 195
R1206 VSS.n766 VSS.n741 195
R1207 VSS.n766 VSS.n765 195
R1208 VSS.n155 VSS.n150 195
R1209 VSS.n1251 VSS.n1250 195
R1210 VSS.n1252 VSS.n1251 195
R1211 VSS.n332 VSS.n331 195
R1212 VSS.n847 VSS.n846 195
R1213 VSS.n1440 VSS.n1439 195
R1214 VSS.n1439 VSS.n1438 195
R1215 VSS.n606 VSS.n603 195
R1216 VSS.n1013 VSS.n1012 194.941
R1217 VSS.n1023 VSS.n1019 194.941
R1218 VSS.n1186 VSS.n1185 194.941
R1219 VSS.n1264 VSS.n1263 194.941
R1220 VSS.n1019 VSS.n492 194.489
R1221 VSS.n1263 VSS.n231 194.489
R1222 VSS.n1013 VSS.n441 189.964
R1223 VSS.n1185 VSS.n201 189.964
R1224 VSS.n664 VSS.n630 181.212
R1225 VSS.n638 VSS.n636 175.543
R1226 VSS.n1122 VSS.n380 175.543
R1227 VSS.n448 VSS.n447 172.892
R1228 VSS.n670 VSS.n669 172.168
R1229 VSS.n1248 VSS 165.862
R1230 VSS.n816 VSS.n736 163.032
R1231 VSS.n777 VSS.n738 163.032
R1232 VSS.n772 VSS.n739 163.032
R1233 VSS.n820 VSS.n819 163.032
R1234 VSS.n943 VSS.n942 162.72
R1235 VSS.n254 VSS.n253 151.356
R1236 VSS.n60 VSS.n58 150.798
R1237 VSS.n556 VSS.t235 147.376
R1238 VSS.t169 VSS.n244 147.376
R1239 VSS.t215 VSS.t235 144.576
R1240 VSS.t237 VSS.t169 144.576
R1241 VSS.n301 VSS.n300 142.526
R1242 VSS.n475 VSS.n473 142.526
R1243 VSS.n816 VSS.n815 139.733
R1244 VSS.n777 VSS.n776 139.733
R1245 VSS.n772 VSS.n771 139.733
R1246 VSS.n821 VSS.n820 139.733
R1247 VSS.n1231 VSS.n179 132.096
R1248 VSS.n1233 VSS.n1232 132.096
R1249 VSS.n1234 VSS.n1230 132.096
R1250 VSS.n1235 VSS.n1229 132.096
R1251 VSS.n1236 VSS.n1228 132.096
R1252 VSS.n1239 VSS.n259 132.096
R1253 VSS.n1240 VSS.n258 132.096
R1254 VSS.n1241 VSS.n257 132.096
R1255 VSS.n1242 VSS.n256 132.096
R1256 VSS.n1243 VSS.n255 132.096
R1257 VSS.n1244 VSS.n254 132.096
R1258 VSS.n1156 VSS.n358 132.096
R1259 VSS.n1157 VSS.n357 132.096
R1260 VSS.n1158 VSS.n356 132.096
R1261 VSS.n1159 VSS.n355 132.096
R1262 VSS.n1160 VSS.n354 132.096
R1263 VSS.n759 VSS.n353 132.096
R1264 VSS.n758 VSS.n744 132.096
R1265 VSS.n757 VSS.n745 132.096
R1266 VSS.n756 VSS.n746 132.096
R1267 VSS.n755 VSS.n747 132.096
R1268 VSS.n754 VSS.n748 132.096
R1269 VSS.n958 VSS.n53 132.096
R1270 VSS.n960 VSS.n959 132.096
R1271 VSS.n961 VSS.n957 132.096
R1272 VSS.n962 VSS.n956 132.096
R1273 VSS.n963 VSS.n955 132.096
R1274 VSS.n983 VSS.n966 132.096
R1275 VSS.n982 VSS.n967 132.096
R1276 VSS.n981 VSS.n968 132.096
R1277 VSS.n980 VSS.n969 132.096
R1278 VSS.n979 VSS.n970 132.096
R1279 VSS.n978 VSS.n971 132.096
R1280 VSS.n1411 VSS.n44 132.096
R1281 VSS.n1412 VSS.n43 132.096
R1282 VSS.n1413 VSS.n42 132.096
R1283 VSS.n1414 VSS.n41 132.096
R1284 VSS.n1415 VSS.n40 132.096
R1285 VSS.n1249 VSS.n1248 129.779
R1286 VSS.n1057 VSS.n1056 129.005
R1287 VSS.n1323 VSS.n158 124.475
R1288 VSS.n122 VSS.n115 124.475
R1289 VSS.n1378 VSS.n92 124.475
R1290 VSS.n840 VSS.n717 124.475
R1291 VSS.n340 VSS.n339 124.475
R1292 VSS.n876 VSS.n875 124.475
R1293 VSS VSS.n200 123.603
R1294 VSS.n160 VSS.n151 122.175
R1295 VSS.n1351 VSS.n1350 122.175
R1296 VSS.n782 VSS.n781 122.175
R1297 VSS.n719 VSS.n712 122.175
R1298 VSS.n335 VSS.n322 122.175
R1299 VSS.n874 VSS.n604 122.175
R1300 VSS.n1222 VSS.n1221 121.922
R1301 VSS.n1394 VSS.n1393 121.922
R1302 VSS.n1389 VSS.n75 121.922
R1303 VSS.n1217 VSS.n274 121.922
R1304 VSS.n359 VSS.n358 121.734
R1305 VSS.n1411 VSS.n1410 121.734
R1306 VSS.n1406 VSS.n53 121.734
R1307 VSS.n1306 VSS.n179 121.734
R1308 VSS.n754 VSS.n753 120.623
R1309 VSS.n972 VSS.n971 120.623
R1310 VSS.n550 VSS.n546 120.367
R1311 VSS.n926 VSS.n923 120.055
R1312 VSS.n546 VSS.n545 119.66
R1313 VSS.n499 VSS.n439 119.04
R1314 VSS.n498 VSS.n443 117.001
R1315 VSS.n443 VSS.t182 117.001
R1316 VSS.n678 VSS.n677 117.001
R1317 VSS.n678 VSS.t119 117.001
R1318 VSS.n1055 VSS.n1054 117.001
R1319 VSS.n1054 VSS.t182 117.001
R1320 VSS.n681 VSS.n680 117.001
R1321 VSS.n680 VSS.t119 117.001
R1322 VSS.n1168 VSS.n204 117.001
R1323 VSS.t23 VSS.n204 117.001
R1324 VSS.n1170 VSS.n318 117.001
R1325 VSS.t146 VSS.n318 117.001
R1326 VSS.n1290 VSS.n1289 117.001
R1327 VSS.n1289 VSS.t23 117.001
R1328 VSS.n1149 VSS.n319 117.001
R1329 VSS.t146 VSS.n319 117.001
R1330 VSS.n1021 VSS.n444 117.001
R1331 VSS.n444 VSS.t182 117.001
R1332 VSS.n994 VSS.n993 117.001
R1333 VSS.n993 VSS.t119 117.001
R1334 VSS.n490 VSS.n445 117.001
R1335 VSS.n445 VSS.t182 117.001
R1336 VSS.n1000 VSS.n999 117.001
R1337 VSS.n999 VSS.t119 117.001
R1338 VSS.n1288 VSS.n1287 117.001
R1339 VSS.t23 VSS.n1288 117.001
R1340 VSS.n1208 VSS.n1207 117.001
R1341 VSS.t146 VSS.n1208 117.001
R1342 VSS.n211 VSS.n205 117.001
R1343 VSS.t23 VSS.n205 117.001
R1344 VSS.n345 VSS.n343 117.001
R1345 VSS.t146 VSS.n343 117.001
R1346 VSS.n832 VSS.n831 117.001
R1347 VSS.t240 VSS.n832 117.001
R1348 VSS.n839 VSS.n838 117.001
R1349 VSS.n838 VSS.t203 117.001
R1350 VSS.n834 VSS.n833 117.001
R1351 VSS.n833 VSS.t240 117.001
R1352 VSS.n837 VSS.n836 117.001
R1353 VSS.t203 VSS.n837 117.001
R1354 VSS.n844 VSS.n843 117.001
R1355 VSS.n843 VSS.t211 117.001
R1356 VSS.n733 VSS.n732 117.001
R1357 VSS.n733 VSS.t167 117.001
R1358 VSS.n817 VSS.n734 117.001
R1359 VSS.n734 VSS.t167 117.001
R1360 VSS.n1370 VSS.n1369 117.001
R1361 VSS.t201 VSS.n1370 117.001
R1362 VSS.n1377 VSS.n1376 117.001
R1363 VSS.n1376 VSS.t78 117.001
R1364 VSS.n1372 VSS.n1371 117.001
R1365 VSS.n1371 VSS.t201 117.001
R1366 VSS.n1375 VSS.n1374 117.001
R1367 VSS.t78 VSS.n1375 117.001
R1368 VSS.n1380 VSS.n1379 117.001
R1369 VSS.t165 VSS.n1380 117.001
R1370 VSS.n800 VSS.n799 117.001
R1371 VSS.t16 VSS.n800 117.001
R1372 VSS.n783 VSS.n88 117.001
R1373 VSS.t165 VSS.n88 117.001
R1374 VSS.n802 VSS.n801 117.001
R1375 VSS.n801 VSS.t16 117.001
R1376 VSS.n106 VSS.n105 117.001
R1377 VSS.t69 VSS.n106 117.001
R1378 VSS.n778 VSS.n107 117.001
R1379 VSS.t69 VSS.n107 117.001
R1380 VSS.n1338 VSS.n1337 117.001
R1381 VSS.t129 VSS.n1338 117.001
R1382 VSS.n141 VSS.n123 117.001
R1383 VSS.t171 VSS.n123 117.001
R1384 VSS.n1340 VSS.n1339 117.001
R1385 VSS.n1339 VSS.t129 117.001
R1386 VSS.n133 VSS.n124 117.001
R1387 VSS.t171 VSS.n124 117.001
R1388 VSS.n1355 VSS.n1354 117.001
R1389 VSS.n1354 VSS.t67 117.001
R1390 VSS.n432 VSS.n114 117.001
R1391 VSS.t218 VSS.n432 117.001
R1392 VSS.n1353 VSS.n1352 117.001
R1393 VSS.t67 VSS.n1353 117.001
R1394 VSS.n429 VSS.n428 117.001
R1395 VSS.t218 VSS.n429 117.001
R1396 VSS.n1335 VSS.n130 117.001
R1397 VSS.t204 VSS.n130 117.001
R1398 VSS.n773 VSS.n131 117.001
R1399 VSS.t204 VSS.n131 117.001
R1400 VSS.n1315 VSS.n1314 117.001
R1401 VSS.t90 VSS.n1315 117.001
R1402 VSS.n1322 VSS.n1321 117.001
R1403 VSS.n1321 VSS.t84 117.001
R1404 VSS.n1317 VSS.n1316 117.001
R1405 VSS.n1316 VSS.t90 117.001
R1406 VSS.n1320 VSS.n1319 117.001
R1407 VSS.t84 VSS.n1320 117.001
R1408 VSS.n1325 VSS.n1324 117.001
R1409 VSS.t206 VSS.n1325 117.001
R1410 VSS.n1333 VSS.n1332 117.001
R1411 VSS.n1332 VSS.t49 117.001
R1412 VSS.n1327 VSS.n1326 117.001
R1413 VSS.n1326 VSS.t206 117.001
R1414 VSS.n1331 VSS.n1330 117.001
R1415 VSS.t49 VSS.n1331 117.001
R1416 VSS.n171 VSS.n170 117.001
R1417 VSS.t135 VSS.n171 117.001
R1418 VSS.n1247 VSS.n172 117.001
R1419 VSS.t135 VSS.n172 117.001
R1420 VSS.n242 VSS.n241 117.001
R1421 VSS.n241 VSS.t115 117.001
R1422 VSS.n342 VSS.n341 117.001
R1423 VSS.t122 VSS.n342 117.001
R1424 VSS.n1256 VSS.n1255 117.001
R1425 VSS.n1255 VSS.t115 117.001
R1426 VSS.n320 VSS.n239 117.001
R1427 VSS.t122 VSS.n320 117.001
R1428 VSS.n323 VSS.n192 117.001
R1429 VSS.t133 VSS.n323 117.001
R1430 VSS.n1300 VSS.n1299 117.001
R1431 VSS.t73 VSS.n1300 117.001
R1432 VSS.n337 VSS.n336 117.001
R1433 VSS.n337 VSS.t133 117.001
R1434 VSS.n325 VSS.n188 117.001
R1435 VSS.t73 VSS.n188 117.001
R1436 VSS.n695 VSS.n694 117.001
R1437 VSS.t213 VSS.n695 117.001
R1438 VSS.n842 VSS.n841 117.001
R1439 VSS.t211 VSS.n842 117.001
R1440 VSS.n715 VSS.n697 117.001
R1441 VSS.t175 VSS.n697 117.001
R1442 VSS.n706 VSS.n698 117.001
R1443 VSS.t175 VSS.n698 117.001
R1444 VSS.n859 VSS.n0 117.001
R1445 VSS.n859 VSS.t213 117.001
R1446 VSS.n867 VSS.n866 117.001
R1447 VSS.n866 VSS.t96 117.001
R1448 VSS.n619 VSS.n613 117.001
R1449 VSS.t239 VSS.n613 117.001
R1450 VSS.n865 VSS.n864 117.001
R1451 VSS.t96 VSS.n865 117.001
R1452 VSS.n612 VSS.n611 117.001
R1453 VSS.t239 VSS.n612 117.001
R1454 VSS.n880 VSS.n879 117.001
R1455 VSS.n879 VSS.t82 117.001
R1456 VSS.n878 VSS.n877 117.001
R1457 VSS.t82 VSS.n878 117.001
R1458 VSS.n598 VSS.n596 117.001
R1459 VSS.n598 VSS.t188 117.001
R1460 VSS.n891 VSS.n890 117.001
R1461 VSS.t109 VSS.n891 117.001
R1462 VSS.n600 VSS.n592 117.001
R1463 VSS.t109 VSS.n592 117.001
R1464 VSS.n884 VSS.n883 117.001
R1465 VSS.n884 VSS.t188 117.001
R1466 VSS.n294 VSS.n292 116.254
R1467 VSS.n1038 VSS.n1037 116.254
R1468 VSS.n194 VSS.n144 113.775
R1469 VSS.n1357 VSS.n1356 113.775
R1470 VSS.n786 VSS.n91 113.775
R1471 VSS.n716 VSS.n705 113.775
R1472 VSS.n701 VSS.n610 113.775
R1473 VSS.n943 VSS.n923 113.59
R1474 VSS.n1057 VSS.n440 112.001
R1475 VSS.n629 VSS.n628 111.27
R1476 VSS.n624 VSS.n528 111.27
R1477 VSS.n348 VSS.n347 110.674
R1478 VSS.n513 VSS.n512 110.674
R1479 VSS.n688 VSS.n670 109.183
R1480 VSS.n1056 VSS.n362 109.183
R1481 VSS.n1291 VSS.n200 109.106
R1482 VSS.n438 VSS.n406 108.745
R1483 VSS.n1285 VSS.n1284 108.299
R1484 VSS.n1284 VSS.n1283 108.186
R1485 VSS.n1429 VSS.n22 107.79
R1486 VSS.n948 VSS.n947 107.79
R1487 VSS.n1109 VSS.n1108 107.79
R1488 VSS.n423 VSS.n421 107.79
R1489 VSS.n1096 VSS.n1095 107.621
R1490 VSS.n1298 VSS.n1297 100.677
R1491 VSS.n601 VSS.n1 99.8
R1492 VSS.n1020 VSS.n488 97.9434
R1493 VSS.n502 VSS.n501 97.9434
R1494 VSS.n1286 VSS.n209 97.9434
R1495 VSS.n1167 VSS.n1166 97.9434
R1496 VSS.n1388 VSS.n1387 97.5005
R1497 VSS.n1387 VSS.n72 97.5005
R1498 VSS.n511 VSS.n78 97.5005
R1499 VSS.n78 VSS.n72 97.5005
R1500 VSS.n1216 VSS.n1215 97.5005
R1501 VSS.n1215 VSS.n271 97.5005
R1502 VSS.n346 VSS.n277 97.5005
R1503 VSS.n277 VSS.n271 97.5005
R1504 VSS.n82 VSS.n67 97.5005
R1505 VSS.n82 VSS.n72 97.5005
R1506 VSS.n475 VSS.n81 97.5005
R1507 VSS.n81 VSS.n72 97.5005
R1508 VSS.n281 VSS.n266 97.5005
R1509 VSS.n281 VSS.n271 97.5005
R1510 VSS.n301 VSS.n280 97.5005
R1511 VSS.n280 VSS.n271 97.5005
R1512 VSS.t62 VSS.t102 89.969
R1513 VSS.t184 VSS.t112 89.969
R1514 VSS.t164 VSS.t100 89.969
R1515 VSS.t100 VSS.t170 89.969
R1516 VSS.t170 VSS.t158 89.969
R1517 VSS.t158 VSS.t65 89.969
R1518 VSS.t65 VSS.t44 89.969
R1519 VSS.t44 VSS.t35 89.969
R1520 VSS.t35 VSS.t5 89.969
R1521 VSS.t5 VSS.t85 89.969
R1522 VSS.t85 VSS.t178 89.969
R1523 VSS.t178 VSS.t98 89.969
R1524 VSS.t98 VSS.t14 89.969
R1525 VSS.t14 VSS.t61 89.969
R1526 VSS.t61 VSS.t64 89.969
R1527 VSS.t64 VSS.t131 89.969
R1528 VSS.t131 VSS.t152 89.969
R1529 VSS.t152 VSS.t7 89.969
R1530 VSS.t7 VSS.t59 89.969
R1531 VSS.t59 VSS.t94 89.969
R1532 VSS.t94 VSS.t142 89.969
R1533 VSS.t142 VSS.t107 89.969
R1534 VSS.t107 VSS.t180 89.969
R1535 VSS.t180 VSS.t24 89.969
R1536 VSS.t24 VSS.t217 89.969
R1537 VSS.t217 VSS.t38 89.969
R1538 VSS.t38 VSS.t114 89.969
R1539 VSS.t114 VSS.t137 89.969
R1540 VSS.t137 VSS.t177 89.969
R1541 VSS.t177 VSS.t63 89.969
R1542 VSS.t63 VSS.t62 89.969
R1543 VSS.t27 VSS.t40 89.969
R1544 VSS.t40 VSS.t157 89.969
R1545 VSS.t157 VSS.t150 89.969
R1546 VSS.t150 VSS.t8 89.969
R1547 VSS.t8 VSS.t143 89.969
R1548 VSS.t143 VSS.t43 89.969
R1549 VSS.t43 VSS.t13 89.969
R1550 VSS.t13 VSS.t126 89.969
R1551 VSS.t126 VSS.t145 89.969
R1552 VSS.t145 VSS.t4 89.969
R1553 VSS.t4 VSS.t104 89.969
R1554 VSS.t104 VSS.t6 89.969
R1555 VSS.t6 VSS.t118 89.969
R1556 VSS.t118 VSS.t160 89.969
R1557 VSS.t160 VSS.t0 89.969
R1558 VSS.t0 VSS.t91 89.969
R1559 VSS.t91 VSS.t174 89.969
R1560 VSS.t174 VSS.t141 89.969
R1561 VSS.t141 VSS.t79 89.969
R1562 VSS.t79 VSS.t39 89.969
R1563 VSS.t39 VSS.t77 89.969
R1564 VSS.t77 VSS.t60 89.969
R1565 VSS.t60 VSS.t116 89.969
R1566 VSS.t116 VSS.t30 89.969
R1567 VSS.t30 VSS.t184 89.969
R1568 VSS.t112 VSS.t57 89.969
R1569 VSS.t57 VSS.t42 89.969
R1570 VSS.t42 VSS.t29 89.969
R1571 VSS.t29 VSS.t51 89.969
R1572 VSS.t51 VSS.t199 89.969
R1573 VSS.n1123 VSS.n377 89.9662
R1574 VSS.n644 VSS.n640 89.9662
R1575 VSS.n1124 VSS.n1122 88.2291
R1576 VSS.n639 VSS.n638 88.2291
R1577 VSS.n830 VSS.n829 87.2389
R1578 VSS.n1368 VSS.n1367 87.2389
R1579 VSS.n1336 VSS.n132 87.2389
R1580 VSS.n1313 VSS.n1312 87.2389
R1581 VSS.n863 VSS.n862 87.2389
R1582 VSS.n1206 VSS.n1205 85.3465
R1583 VSS.n996 VSS.n995 85.3465
R1584 VSS.n675 VSS.n76 85.3465
R1585 VSS.n1144 VSS.n275 85.3465
R1586 VSS.n1245 VSS.n1244 84.1782
R1587 VSS.n552 VSS.n550 82.0392
R1588 VSS.t132 VSS.n893 81.126
R1589 VSS.n554 VSS.n545 80.7449
R1590 VSS.t201 VSS.n103 80.5207
R1591 VSS.n1441 VSS.n1 79.8295
R1592 VSS.n1049 VSS.n1048 78.6291
R1593 VSS.n1282 VSS.n1281 78.6291
R1594 VSS.n828 VSS.n726 77.6035
R1595 VSS.n1366 VSS.n100 77.6035
R1596 VSS.n1342 VSS.n1341 77.6035
R1597 VSS.n1311 VSS.n166 77.6035
R1598 VSS.n861 VSS.n2 77.6035
R1599 VSS.n629 VSS.n21 76.8005
R1600 VSS.n624 VSS.n527 76.8005
R1601 VSS.n543 VSS.t215 72.2878
R1602 VSS.n543 VSS.t237 72.2878
R1603 VSS.n1188 VSS.n274 72.1925
R1604 VSS.n1190 VSS.n1189 72.1925
R1605 VSS.n1191 VSS.n1164 72.1925
R1606 VSS.n1192 VSS.n1163 72.1925
R1607 VSS.n1193 VSS.n1162 72.1925
R1608 VSS.n1197 VSS.n1196 72.1925
R1609 VSS.n1198 VSS.n352 72.1925
R1610 VSS.n1199 VSS.n351 72.1925
R1611 VSS.n1200 VSS.n350 72.1925
R1612 VSS.n1201 VSS.n349 72.1925
R1613 VSS.n1202 VSS.n348 72.1925
R1614 VSS.n1222 VSS.n228 72.1925
R1615 VSS.n1223 VSS.n227 72.1925
R1616 VSS.n1224 VSS.n265 72.1925
R1617 VSS.n1225 VSS.n264 72.1925
R1618 VSS.n1226 VSS.n263 72.1925
R1619 VSS.n295 VSS.n282 72.1925
R1620 VSS.n296 VSS.n285 72.1925
R1621 VSS.n297 VSS.n287 72.1925
R1622 VSS.n298 VSS.n289 72.1925
R1623 VSS.n299 VSS.n291 72.1925
R1624 VSS.n300 VSS.n293 72.1925
R1625 VSS.n1394 VSS.n66 72.1925
R1626 VSS.n1395 VSS.n65 72.1925
R1627 VSS.n1396 VSS.n64 72.1925
R1628 VSS.n1397 VSS.n63 72.1925
R1629 VSS.n1398 VSS.n62 72.1925
R1630 VSS.n468 VSS.n83 72.1925
R1631 VSS.n481 VSS.n469 72.1925
R1632 VSS.n480 VSS.n470 72.1925
R1633 VSS.n479 VSS.n471 72.1925
R1634 VSS.n478 VSS.n472 72.1925
R1635 VSS.n477 VSS.n473 72.1925
R1636 VSS.n503 VSS.n75 72.1925
R1637 VSS.n518 VSS.n505 72.1925
R1638 VSS.n519 VSS.n507 72.1925
R1639 VSS.n520 VSS.n509 72.1925
R1640 VSS.n521 VSS.n510 72.1925
R1641 VSS.n986 VSS.n985 72.1925
R1642 VSS.n987 VSS.n517 72.1925
R1643 VSS.n988 VSS.n516 72.1925
R1644 VSS.n989 VSS.n515 72.1925
R1645 VSS.n990 VSS.n514 72.1925
R1646 VSS.n991 VSS.n513 72.1925
R1647 VSS.n895 VSS.t132 69.976
R1648 VSS.n915 VSS.t199 69.976
R1649 VSS.n664 VSS.n663 67.742
R1650 VSS.n688 VSS.n687 66.8449
R1651 VSS.n687 VSS.n686 66.8449
R1652 VSS.n1141 VSS.n362 66.8449
R1653 VSS.n1142 VSS.n1141 66.8449
R1654 VSS.n1390 VSS.n1389 65.0005
R1655 VSS.n1391 VSS.n1390 65.0005
R1656 VSS.n683 VSS.n71 65.0005
R1657 VSS.n1391 VSS.n71 65.0005
R1658 VSS.n1218 VSS.n1217 65.0005
R1659 VSS.n1219 VSS.n1218 65.0005
R1660 VSS.n1151 VSS.n270 65.0005
R1661 VSS.n1219 VSS.n270 65.0005
R1662 VSS.n1393 VSS.n1392 65.0005
R1663 VSS.n1392 VSS.n1391 65.0005
R1664 VSS.n512 VSS.n70 65.0005
R1665 VSS.n1391 VSS.n70 65.0005
R1666 VSS.n1221 VSS.n1220 65.0005
R1667 VSS.n1220 VSS.n1219 65.0005
R1668 VSS.n347 VSS.n269 65.0005
R1669 VSS.n1219 VSS.n269 65.0005
R1670 VSS.n1078 VSS.n1076 64.0005
R1671 VSS.n1076 VSS.n1074 64.0005
R1672 VSS.n1074 VSS.n1072 64.0005
R1673 VSS.n1072 VSS.n1070 64.0005
R1674 VSS.n1070 VSS.n410 64.0005
R1675 VSS.n1101 VSS.n1100 64.0005
R1676 VSS.n1100 VSS.n1099 64.0005
R1677 VSS.n1099 VSS.n1098 64.0005
R1678 VSS.n1098 VSS.n1097 64.0005
R1679 VSS.n665 VSS.n664 63.8619
R1680 VSS.n665 VSS.n629 63.756
R1681 VSS.n669 VSS.n624 63.756
R1682 VSS.n302 VSS.n301 63.3268
R1683 VSS.n476 VSS.n475 63.3268
R1684 VSS.n1204 VSS.n1203 60.2167
R1685 VSS.n997 VSS.n992 60.2167
R1686 VSS.n977 VSS.n976 59.7818
R1687 VSS.n751 VSS.n750 59.7818
R1688 VSS.t185 VSS.t36 59.2846
R1689 VSS.t37 VSS.n768 59.2846
R1690 VSS.n673 VSS.n54 58.8258
R1691 VSS.n975 VSS.n974 58.8258
R1692 VSS.n749 VSS.n180 58.8258
R1693 VSS.n1155 VSS.n1154 58.8258
R1694 VSS.n690 VSS.n32 58.1547
R1695 VSS.n1428 VSS.n23 58.1547
R1696 VSS.n425 VSS.n424 58.1547
R1697 VSS.n1061 VSS.n364 58.1547
R1698 VSS.n607 VSS.t227 57.8099
R1699 VSS.n902 VSS.n901 57.6785
R1700 VSS.t22 VSS.t179 57.5149
R1701 VSS.n682 VSS.n676 57.2498
R1702 VSS.n1150 VSS.n1148 57.2498
R1703 VSS.n1245 VSS.n253 57.0391
R1704 VSS.n644 VSS.n643 56.8991
R1705 VSS.n1127 VSS.n377 56.8991
R1706 VSS.n642 VSS.n641 56.5484
R1707 VSS.n671 VSS.n33 56.5484
R1708 VSS.n367 VSS.n366 56.5484
R1709 VSS.n1129 VSS.n1128 56.5484
R1710 VSS.n638 VSS.n637 56.5458
R1711 VSS.n1122 VSS.n381 56.5458
R1712 VSS.n1063 VSS.n148 56.2422
R1713 VSS.n1361 VSS.n109 56.2422
R1714 VSS.n796 VSS.n737 56.2422
R1715 VSS.n251 VSS.n250 56.2422
R1716 VSS.n854 VSS.n700 56.2422
R1717 VSS.n601 VSS.n597 56.2422
R1718 VSS.n684 VSS.n674 56.1978
R1719 VSS.n1153 VSS.n1152 56.1978
R1720 VSS.n826 VSS.t209 55.7452
R1721 VSS.n1012 VSS.n1011 55.4025
R1722 VSS.n1024 VSS.n1023 55.4025
R1723 VSS.n1187 VSS.n1186 55.4025
R1724 VSS.n1265 VSS.n1264 55.4025
R1725 VSS.n125 VSS.t48 54.8604
R1726 VSS.n1334 VSS.n143 54.5229
R1727 VSS.n113 VSS.n108 54.5229
R1728 VSS.n798 VSS.n797 54.5229
R1729 VSS.n247 VSS.n191 54.5229
R1730 VSS.n855 VSS.n699 54.5229
R1731 VSS.n889 VSS.n888 54.5229
R1732 VSS.n1130 VSS.n1129 54.2902
R1733 VSS.n1422 VSS.n33 54.2902
R1734 VSS.n641 VSS.n24 54.2902
R1735 VSS.n1136 VSS.n367 54.2902
R1736 VSS.n1067 VSS.n1066 54.2705
R1737 VSS.n689 VSS.n688 53.8306
R1738 VSS.n686 VSS.n672 53.8306
R1739 VSS.n1060 VSS.n362 53.8306
R1740 VSS.n1142 VSS.n361 53.8306
R1741 VSS.n625 VSS.t144 53.6806
R1742 VSS.n1385 VSS.t192 53.6806
R1743 VSS.n1105 VSS.t172 53.6806
R1744 VSS.n1090 VSS.t208 53.6806
R1745 VSS.n1213 VSS.t41 53.6806
R1746 VSS.t122 VSS.n233 53.6806
R1747 VSS.n235 VSS.t163 53.6806
R1748 VSS.t230 VSS.n714 53.3857
R1749 VSS.n424 VSS.n375 53.2419
R1750 VSS.n1423 VSS.n32 53.2419
R1751 VSS.n1428 VSS.n1427 53.2419
R1752 VSS.n1137 VSS.n364 53.2419
R1753 VSS.t95 VSS.t21 52.2059
R1754 VSS.n1438 VSS.n1437 52.2059
R1755 VSS.t211 VSS.t229 51.9109
R1756 VSS.n1442 VSS.n0 51.8555
R1757 VSS.n601 VSS.n600 51.6506
R1758 VSS.n902 VSS.n577 51.5907
R1759 VSS.n818 VSS.n817 51.3352
R1760 VSS.n779 VSS.n778 51.3352
R1761 VSS.n774 VSS.n773 51.3352
R1762 VSS.n1273 VSS.t115 51.321
R1763 VSS.n580 VSS.n576 51.2781
R1764 VSS.t84 VSS.t32 50.7312
R1765 VSS.n573 VSS.n571 50.5799
R1766 VSS.n909 VSS.n908 50.5799
R1767 VSS.t148 VSS.t20 50.4362
R1768 VSS.n1247 VSS.n1246 50.2573
R1769 VSS.n248 VSS.t127 50.1413
R1770 VSS.n583 VSS.n573 49.9087
R1771 VSS.n908 VSS.n572 49.649
R1772 VSS.n578 VSS.n576 49.5714
R1773 VSS.n566 VSS.n565 49.1835
R1774 VSS.n563 VSS.n561 49.1835
R1775 VSS.n922 VSS.n921 49.0284
R1776 VSS.n492 VSS.n450 49.0025
R1777 VSS.n231 VSS.n212 49.0025
R1778 VSS.t78 VSS.n96 48.6665
R1779 VSS.n1015 VSS.t173 48.3716
R1780 VSS.t149 VSS.n1003 47.1918
R1781 VSS.n752 VSS.n751 47.1776
R1782 VSS.n977 VSS.n973 47.1776
R1783 VSS.t11 VSS.t66 46.8969
R1784 VSS.t96 VSS.n693 46.8969
R1785 VSS.n1402 VSS.t75 46.8969
R1786 VSS.t240 VSS.t101 46.307
R1787 VSS.t161 VSS.n858 45.7171
R1788 VSS.n848 VSS.t128 45.7171
R1789 VSS.t12 VSS.t92 45.1272
R1790 VSS.t242 VSS.t243 45.1272
R1791 VSS.n1405 VSS.n1404 45.0005
R1792 VSS.n1404 VSS.n50 45.0005
R1793 VSS.n973 VSS.n56 45.0005
R1794 VSS.n56 VSS.n50 45.0005
R1795 VSS.n743 VSS.n360 45.0005
R1796 VSS.n743 VSS.n175 45.0005
R1797 VSS.n752 VSS.n742 45.0005
R1798 VSS.n742 VSS.n175 45.0005
R1799 VSS.n59 VSS.n45 45.0005
R1800 VSS.n59 VSS.n50 45.0005
R1801 VSS.n58 VSS.n50 45.0005
R1802 VSS.n1305 VSS.n1304 45.0005
R1803 VSS.n1304 VSS.n175 45.0005
R1804 VSS.n253 VSS.n182 45.0005
R1805 VSS.n182 VSS.n175 45.0005
R1806 VSS.n905 VSS.t102 44.9848
R1807 VSS.n905 VSS.t27 44.9848
R1808 VSS.n812 VSS.t9 44.8322
R1809 VSS.n464 VSS.n463 44.8005
R1810 VSS.n305 VSS.n304 44.8005
R1811 VSS.n1348 VSS.t210 44.5373
R1812 VSS.n958 VSS.n54 44.4933
R1813 VSS.n974 VSS.n44 44.4933
R1814 VSS.n1231 VSS.n180 44.4933
R1815 VSS.n1156 VSS.n1155 44.4933
R1816 VSS.t246 VSS.t81 43.3575
R1817 VSS.n886 VSS.t33 43.3575
R1818 VSS.n1209 VSS.t139 43.3575
R1819 VSS.n793 VSS.n791 43.3575
R1820 VSS.n1419 VSS.n37 43.0626
R1821 VSS.n1133 VSS.n168 43.0626
R1822 VSS.n767 VSS.t80 42.7676
R1823 VSS.n439 VSS.n438 42.3336
R1824 VSS.n1265 VSS.n209 42.2405
R1825 VSS.n1267 VSS.n1266 42.2405
R1826 VSS.n1268 VSS.n226 42.2405
R1827 VSS.n1269 VSS.n225 42.2405
R1828 VSS.n1270 VSS.n224 42.2405
R1829 VSS.n310 VSS.n223 42.2405
R1830 VSS.n309 VSS.n284 42.2405
R1831 VSS.n308 VSS.n286 42.2405
R1832 VSS.n307 VSS.n288 42.2405
R1833 VSS.n306 VSS.n290 42.2405
R1834 VSS.n305 VSS.n292 42.2405
R1835 VSS.n1187 VSS.n1166 42.2405
R1836 VSS.n1175 VSS.n1165 42.2405
R1837 VSS.n1177 VSS.n1176 42.2405
R1838 VSS.n1178 VSS.n1174 42.2405
R1839 VSS.n1179 VSS.n1173 42.2405
R1840 VSS.n1276 VSS.n217 42.2405
R1841 VSS.n1277 VSS.n216 42.2405
R1842 VSS.n1278 VSS.n215 42.2405
R1843 VSS.n1279 VSS.n214 42.2405
R1844 VSS.n1280 VSS.n213 42.2405
R1845 VSS.n1188 VSS.n1187 42.2405
R1846 VSS.n1189 VSS.n1165 42.2405
R1847 VSS.n1177 VSS.n1164 42.2405
R1848 VSS.n1178 VSS.n1163 42.2405
R1849 VSS.n1179 VSS.n1162 42.2405
R1850 VSS.n1197 VSS.n217 42.2405
R1851 VSS.n1198 VSS.n216 42.2405
R1852 VSS.n1199 VSS.n215 42.2405
R1853 VSS.n1200 VSS.n214 42.2405
R1854 VSS.n1201 VSS.n213 42.2405
R1855 VSS.n1265 VSS.n228 42.2405
R1856 VSS.n1266 VSS.n227 42.2405
R1857 VSS.n265 VSS.n226 42.2405
R1858 VSS.n264 VSS.n225 42.2405
R1859 VSS.n263 VSS.n224 42.2405
R1860 VSS.n310 VSS.n282 42.2405
R1861 VSS.n309 VSS.n285 42.2405
R1862 VSS.n308 VSS.n287 42.2405
R1863 VSS.n307 VSS.n289 42.2405
R1864 VSS.n306 VSS.n291 42.2405
R1865 VSS.n305 VSS.n293 42.2405
R1866 VSS.n1024 VSS.n488 42.2405
R1867 VSS.n1025 VSS.n487 42.2405
R1868 VSS.n1026 VSS.n486 42.2405
R1869 VSS.n1027 VSS.n485 42.2405
R1870 VSS.n1028 VSS.n484 42.2405
R1871 VSS.n1032 VSS.n1030 42.2405
R1872 VSS.n1033 VSS.n482 42.2405
R1873 VSS.n1034 VSS.n467 42.2405
R1874 VSS.n1035 VSS.n466 42.2405
R1875 VSS.n1036 VSS.n465 42.2405
R1876 VSS.n1037 VSS.n464 42.2405
R1877 VSS.n1011 VSS.n502 42.2405
R1878 VSS.n1010 VSS.n504 42.2405
R1879 VSS.n1009 VSS.n506 42.2405
R1880 VSS.n1008 VSS.n508 42.2405
R1881 VSS.n1007 VSS.n456 42.2405
R1882 VSS.n1043 VSS.n455 42.2405
R1883 VSS.n1044 VSS.n454 42.2405
R1884 VSS.n1045 VSS.n453 42.2405
R1885 VSS.n1046 VSS.n452 42.2405
R1886 VSS.n1047 VSS.n451 42.2405
R1887 VSS.n1048 VSS.n450 42.2405
R1888 VSS.n1011 VSS.n503 42.2405
R1889 VSS.n1010 VSS.n505 42.2405
R1890 VSS.n1009 VSS.n507 42.2405
R1891 VSS.n1008 VSS.n509 42.2405
R1892 VSS.n1007 VSS.n510 42.2405
R1893 VSS.n986 VSS.n455 42.2405
R1894 VSS.n987 VSS.n454 42.2405
R1895 VSS.n988 VSS.n453 42.2405
R1896 VSS.n989 VSS.n452 42.2405
R1897 VSS.n990 VSS.n451 42.2405
R1898 VSS.n991 VSS.n450 42.2405
R1899 VSS.n1024 VSS.n66 42.2405
R1900 VSS.n1025 VSS.n65 42.2405
R1901 VSS.n1026 VSS.n64 42.2405
R1902 VSS.n1027 VSS.n63 42.2405
R1903 VSS.n1028 VSS.n62 42.2405
R1904 VSS.n1030 VSS.n83 42.2405
R1905 VSS.n482 VSS.n481 42.2405
R1906 VSS.n480 VSS.n467 42.2405
R1907 VSS.n479 VSS.n466 42.2405
R1908 VSS.n478 VSS.n465 42.2405
R1909 VSS.n477 VSS.n464 42.2405
R1910 VSS.n1281 VSS.n212 42.2405
R1911 VSS.n1202 VSS.n212 42.2405
R1912 VSS.n1335 VSS.n1334 41.4931
R1913 VSS.n113 VSS.n105 41.4931
R1914 VSS.n798 VSS.n732 41.4931
R1915 VSS.n699 VSS.n694 41.4931
R1916 VSS.n890 VSS.n889 41.4931
R1917 VSS.t111 VSS.t25 39.8182
R1918 VSS.t222 VSS.t236 39.8182
R1919 VSS.n1062 VSS.t86 39.8182
R1920 VSS.n641 VSS.n20 39.2772
R1921 VSS.n950 VSS.n33 39.2772
R1922 VSS.n404 VSS.n367 39.2772
R1923 VSS.n1129 VSS.n376 39.2772
R1924 VSS.n978 VSS.n977 38.8101
R1925 VSS.n751 VSS.n748 38.8101
R1926 VSS.n686 VSS.n685 38.6193
R1927 VSS.n685 VSS.n684 38.6193
R1928 VSS.n1143 VSS.n1142 38.6193
R1929 VSS.n1152 VSS.n1143 38.6193
R1930 VSS.n729 VSS.n722 38.3434
R1931 VSS.t49 VSS.t89 38.3434
R1932 VSS.n763 VSS.n169 38.3434
R1933 VSS.n1336 VSS.n1335 38.2856
R1934 VSS.n1368 VSS.n105 38.2856
R1935 VSS.n830 VSS.n732 38.2856
R1936 VSS.n863 VSS.n694 38.2856
R1937 VSS.t56 VSS.t186 38.0485
R1938 VSS.t3 VSS.t197 38.0485
R1939 VSS.t46 VSS.n1363 37.7536
R1940 VSS.n434 VSS.t138 37.7536
R1941 VSS.n330 VSS.n328 37.7536
R1942 VSS.n1250 VSS.n240 37.7148
R1943 VSS.t213 VSS.t125 37.1637
R1944 VSS.n1155 VSS.n360 37.1061
R1945 VSS.n974 VSS.n45 37.1061
R1946 VSS.n1405 VSS.n54 37.1061
R1947 VSS.n1305 VSS.n180 37.1061
R1948 VSS.n304 VSS.n294 37.0531
R1949 VSS.n303 VSS.n302 37.0531
R1950 VSS.n304 VSS.n303 37.0531
R1951 VSS.n1038 VSS.n463 37.0531
R1952 VSS.n476 VSS.n474 37.0531
R1953 VSS.n474 VSS.n463 37.0531
R1954 VSS.n500 VSS.n499 36.8115
R1955 VSS.n60 VSS.n39 36.6792
R1956 VSS.n669 VSS.n668 36.563
R1957 VSS.n668 VSS.n667 36.563
R1958 VSS.n691 VSS.n690 36.563
R1959 VSS.n693 VSS.n691 36.563
R1960 VSS.n689 VSS.n30 36.563
R1961 VSS.n30 VSS.n5 36.563
R1962 VSS.n672 VSS.n31 36.563
R1963 VSS.n37 VSS.n31 36.563
R1964 VSS.n1059 VSS.n1058 36.563
R1965 VSS.n1059 VSS.n104 36.563
R1966 VSS.n1091 VSS.n1061 36.563
R1967 VSS.n1091 VSS.n1090 36.563
R1968 VSS.n1060 VSS.n363 36.563
R1969 VSS.n1067 VSS.n363 36.563
R1970 VSS.n1139 VSS.n361 36.563
R1971 VSS.n1139 VSS.n168 36.563
R1972 VSS.n666 VSS.n665 36.563
R1973 VSS.n667 VSS.n666 36.563
R1974 VSS.n621 VSS.n23 36.563
R1975 VSS.n693 VSS.n621 36.563
R1976 VSS.n637 VSS.n25 36.563
R1977 VSS.n25 VSS.n5 36.563
R1978 VSS.n643 VSS.n26 36.563
R1979 VSS.n37 VSS.n26 36.563
R1980 VSS.n422 VSS.n420 36.563
R1981 VSS.n422 VSS.n104 36.563
R1982 VSS.n426 VSS.n425 36.563
R1983 VSS.n1090 VSS.n426 36.563
R1984 VSS.n381 VSS.n379 36.563
R1985 VSS.n1067 VSS.n379 36.563
R1986 VSS.n1127 VSS.n1126 36.563
R1987 VSS.n1126 VSS.n168 36.563
R1988 VSS.n1324 VSS.n1323 36.4134
R1989 VSS.n1355 VSS.n115 36.4134
R1990 VSS.n1379 VSS.n1378 36.4134
R1991 VSS.n841 VSS.n840 36.4134
R1992 VSS.n877 VSS.n876 36.4134
R1993 VSS.t25 VSS.t202 36.2788
R1994 VSS.t34 VSS.t171 35.9839
R1995 VSS.n1206 VSS.n228 35.8998
R1996 VSS.n995 VSS.n66 35.8998
R1997 VSS.n503 VSS.n76 35.8998
R1998 VSS.n1188 VSS.n275 35.8998
R1999 VSS.n1102 VSS.n1101 35.5205
R2000 VSS.n949 VSS.n948 34.6769
R2001 VSS.n1430 VSS.n1429 34.6769
R2002 VSS.n423 VSS.n419 34.6769
R2003 VSS.n1110 VSS.n1109 34.6769
R2004 VSS.n546 VSS.n542 34.4123
R2005 VSS.n543 VSS.n542 34.4123
R2006 VSS.n553 VSS.n544 34.4123
R2007 VSS.n544 VSS.n543 34.4123
R2008 VSS.n1407 VSS.n1406 34.4123
R2009 VSS.n1408 VSS.n1407 34.4123
R2010 VSS.n671 VSS.n51 34.4123
R2011 VSS.n722 VSS.n51 34.4123
R2012 VSS.n674 VSS.n52 34.4123
R2013 VSS.n789 VSS.n52 34.4123
R2014 VSS.n685 VSS.n49 34.4123
R2015 VSS.n1408 VSS.n49 34.4123
R2016 VSS.n359 VSS.n176 34.4123
R2017 VSS.n1308 VSS.n176 34.4123
R2018 VSS.n366 VSS.n365 34.4123
R2019 VSS.n365 VSS.n169 34.4123
R2020 VSS.n1153 VSS.n186 34.4123
R2021 VSS.n1301 VSS.n186 34.4123
R2022 VSS.n1143 VSS.n174 34.4123
R2023 VSS.n1308 VSS.n174 34.4123
R2024 VSS.n679 VSS.n676 34.4123
R2025 VSS.n679 VSS.n86 34.4123
R2026 VSS.n1014 VSS.n1013 34.4123
R2027 VSS.n1017 VSS.n1014 34.4123
R2028 VSS.n1053 VSS.n440 34.4123
R2029 VSS.n1053 VSS.n1052 34.4123
R2030 VSS.n1148 VSS.n1147 34.4123
R2031 VSS.n1147 VSS.n1146 34.4123
R2032 VSS.n1185 VSS.n234 34.4123
R2033 VSS.n1261 VSS.n234 34.4123
R2034 VSS.n203 VSS.n200 34.4123
R2035 VSS.n220 VSS.n203 34.4123
R2036 VSS.n1410 VSS.n1409 34.4123
R2037 VSS.n1409 VSS.n1408 34.4123
R2038 VSS.n642 VSS.n46 34.4123
R2039 VSS.n722 VSS.n46 34.4123
R2040 VSS.n976 VSS.n47 34.4123
R2041 VSS.n789 VSS.n47 34.4123
R2042 VSS.n972 VSS.n48 34.4123
R2043 VSS.n1408 VSS.n48 34.4123
R2044 VSS.n1307 VSS.n1306 34.4123
R2045 VSS.n1308 VSS.n1307 34.4123
R2046 VSS.n1128 VSS.n177 34.4123
R2047 VSS.n177 VSS.n169 34.4123
R2048 VSS.n750 VSS.n178 34.4123
R2049 VSS.n1301 VSS.n178 34.4123
R2050 VSS.n753 VSS.n173 34.4123
R2051 VSS.n1308 VSS.n173 34.4123
R2052 VSS.n998 VSS.n997 34.4123
R2053 VSS.n998 VSS.n86 34.4123
R2054 VSS.n1019 VSS.n1018 34.4123
R2055 VSS.n1018 VSS.n1017 34.4123
R2056 VSS.n1051 VSS.n1050 34.4123
R2057 VSS.n1052 VSS.n1051 34.4123
R2058 VSS.n1204 VSS.n344 34.4123
R2059 VSS.n1146 VSS.n344 34.4123
R2060 VSS.n1263 VSS.n1262 34.4123
R2061 VSS.n1262 VSS.n1261 34.4123
R2062 VSS.n1284 VSS.n207 34.4123
R2063 VSS.n220 VSS.n207 34.4123
R2064 VSS.n1334 VSS.n1333 33.8211
R2065 VSS.n114 VSS.n113 33.8211
R2066 VSS.n799 VSS.n798 33.8211
R2067 VSS.n715 VSS.n699 33.8211
R2068 VSS.n889 VSS.n596 33.8211
R2069 VSS.n1333 VSS.n144 33.6319
R2070 VSS.n1356 VSS.n114 33.6319
R2071 VSS.n799 VSS.n91 33.6319
R2072 VSS.n716 VSS.n715 33.6319
R2073 VSS.n610 VSS.n596 33.6319
R2074 VSS.t113 VSS.n531 33.6243
R2075 VSS.n1093 VSS.t183 33.6243
R2076 VSS.n1324 VSS.n144 33.5064
R2077 VSS.n1356 VSS.n1355 33.5064
R2078 VSS.n1379 VSS.n91 33.5064
R2079 VSS.n841 VSS.n716 33.5064
R2080 VSS.n877 VSS.n610 33.5064
R2081 VSS.n645 VSS.n644 33.2279
R2082 VSS.n382 VSS.n377 33.2279
R2083 VSS.n790 VSS.n789 33.0344
R2084 VSS.n1309 VSS.t71 33.0344
R2085 VSS.n328 VSS.n187 33.0344
R2086 VSS.n1146 VSS.n1145 33.0344
R2087 VSS.t202 VSS.t246 32.7395
R2088 VSS.t244 VSS.t46 32.7395
R2089 VSS.n673 VSS.n73 32.5005
R2090 VSS.n790 VSS.n73 32.5005
R2091 VSS.n675 VSS.n74 32.5005
R2092 VSS.n80 VSS.n74 32.5005
R2093 VSS.n1154 VSS.n272 32.5005
R2094 VSS.n272 VSS.n187 32.5005
R2095 VSS.n1144 VSS.n273 32.5005
R2096 VSS.n1145 VSS.n273 32.5005
R2097 VSS.n975 VSS.n68 32.5005
R2098 VSS.n790 VSS.n68 32.5005
R2099 VSS.n996 VSS.n69 32.5005
R2100 VSS.n80 VSS.n69 32.5005
R2101 VSS.n749 VSS.n267 32.5005
R2102 VSS.n267 VSS.n187 32.5005
R2103 VSS.n1205 VSS.n268 32.5005
R2104 VSS.n1145 VSS.n268 32.5005
R2105 VSS.t221 VSS.n72 32.4445
R2106 VSS.t195 VSS.n157 32.4445
R2107 VSS.n992 VSS.n991 32.1277
R2108 VSS.n1203 VSS.n1202 32.1277
R2109 VSS.n405 VSS.n403 32.0005
R2110 VSS.n403 VSS.n401 32.0005
R2111 VSS.n401 VSS.n399 32.0005
R2112 VSS.n399 VSS.n397 32.0005
R2113 VSS.n397 VSS.n396 32.0005
R2114 VSS.n396 VSS.n391 32.0005
R2115 VSS.n391 VSS.n389 32.0005
R2116 VSS.n389 VSS.n387 32.0005
R2117 VSS.n387 VSS.n385 32.0005
R2118 VSS.n385 VSS.n383 32.0005
R2119 VSS.n857 VSS.t190 31.2647
R2120 VSS.n901 VSS.n900 31.22
R2121 VSS.n900 VSS.n538 31.22
R2122 VSS.n919 VSS.n918 31.22
R2123 VSS.n920 VSS.n919 31.22
R2124 VSS.t198 VSS.t97 30.9698
R2125 VSS.t31 VSS.t108 30.9698
R2126 VSS.n693 VSS.n692 30.6749
R2127 VSS.n1408 VSS.t58 30.6749
R2128 VSS.t162 VSS.n1308 30.6749
R2129 VSS.n1302 VSS.n1301 30.6749
R2130 VSS.t125 VSS.t233 30.3799
R2131 VSS.t194 VSS.t130 30.3799
R2132 VSS.t165 VSS.t119 30.085
R2133 VSS.t193 VSS.t175 29.79
R2134 VSS.n430 VSS.t18 29.79
R2135 VSS.t133 VSS.n271 29.79
R2136 VSS.n638 VSS.n631 29.4017
R2137 VSS.n1122 VSS.n1121 29.4017
R2138 VSS.n302 VSS.n293 29.3727
R2139 VSS.n477 VSS.n476 29.3727
R2140 VSS.t66 VSS.t111 29.2001
R2141 VSS.t236 VSS.t69 29.2001
R2142 VSS.t218 VSS.t103 29.2001
R2143 VSS.n1425 VSS.t245 28.9052
R2144 VSS.n1391 VSS.t99 28.9052
R2145 VSS.n156 VSS.t151 28.9052
R2146 VSS.n1219 VSS.t241 28.9052
R2147 VSS.t117 VSS.n857 28.6102
R2148 VSS.n1309 VSS.t147 28.6102
R2149 VSS.t223 VSS.t218 28.3153
R2150 VSS.n449 VSS.n448 27.9585
R2151 VSS.n138 VSS.t31 27.4305
R2152 VSS.n191 VSS.n170 27.2784
R2153 VSS.t120 VSS.t135 27.1355
R2154 VSS.n340 VSS.n192 27.1099
R2155 VSS.n1206 VSS.n266 26.9378
R2156 VSS.n995 VSS.n67 26.9378
R2157 VSS.n1388 VSS.n76 26.9378
R2158 VSS.n1216 VSS.n275 26.9378
R2159 VSS.n942 VSS.n941 26.8805
R2160 VSS.n1082 VSS.n1081 26.8805
R2161 VSS.n1133 VSS.n372 26.8406
R2162 VSS.t186 VSS.n871 26.2507
R2163 VSS.t88 VSS.n155 26.2507
R2164 VSS.t45 VSS.n767 26.2507
R2165 VSS.t123 VSS.n184 26.2507
R2166 VSS.n1301 VSS.t73 26.2507
R2167 VSS.n1256 VSS.n240 25.9798
R2168 VSS.n1052 VSS.n96 25.9557
R2169 VSS.n1273 VSS.n220 25.9557
R2170 VSS.n1203 VSS.n346 25.7834
R2171 VSS.n992 VSS.n511 25.7834
R2172 VSS.t105 VSS.t47 25.6608
R2173 VSS.n4 VSS.n1 25.4353
R2174 VSS.t228 VSS.n4 25.4353
R2175 VSS.n724 VSS.n710 25.4353
R2176 VSS.t140 VSS.n710 25.4353
R2177 VSS.n815 VSS.n814 25.4353
R2178 VSS.n814 VSS.t173 25.4353
R2179 VSS.n809 VSS.n98 25.4353
R2180 VSS.n809 VSS.t173 25.4353
R2181 VSS.n776 VSS.n126 25.4353
R2182 VSS.t224 VSS.n126 25.4353
R2183 VSS.n1347 VSS.n121 25.4353
R2184 VSS.t224 VSS.n1347 25.4353
R2185 VSS.n771 VSS.n770 25.4353
R2186 VSS.n770 VSS.t93 25.4353
R2187 VSS.n769 VSS.n164 25.4353
R2188 VSS.t93 VSS.n769 25.4353
R2189 VSS.n1249 VSS.n246 25.4353
R2190 VSS.t139 VSS.n246 25.4353
R2191 VSS.n334 VSS.n245 25.4353
R2192 VSS.t139 VSS.n245 25.4353
R2193 VSS.n821 VSS.n711 25.4353
R2194 VSS.t140 VSS.n711 25.4353
R2195 VSS.n618 VSS.n3 25.4353
R2196 VSS.t228 VSS.n3 25.4353
R2197 VSS.n1319 VSS.n1318 25.4109
R2198 VSS.n1318 VSS.n1317 25.4109
R2199 VSS.n134 VSS.n133 25.4109
R2200 VSS.n1340 VSS.n134 25.4109
R2201 VSS.n1374 VSS.n1373 25.4109
R2202 VSS.n1373 VSS.n1372 25.4109
R2203 VSS.n836 VSS.n835 25.4109
R2204 VSS.n835 VSS.n834 25.4109
R2205 VSS.n1257 VSS.n239 25.4109
R2206 VSS.n1257 VSS.n1256 25.4109
R2207 VSS.n868 VSS.n619 25.4109
R2208 VSS.n868 VSS.n867 25.4109
R2209 VSS.n1299 VSS.n191 25.3496
R2210 VSS.n684 VSS.n683 24.5065
R2211 VSS.n683 VSS.n682 24.5065
R2212 VSS.n1152 VSS.n1151 24.5065
R2213 VSS.n1151 VSS.n1150 24.5065
R2214 VSS.n794 VSS.n790 24.481
R2215 VSS.n1260 VSS.n235 24.481
R2216 VSS.n1381 VSS.n86 24.186
R2217 VSS.t156 VSS.t12 23.8911
R2218 VSS.t55 VSS.t34 23.8911
R2219 VSS.n1209 VSS.n315 23.8911
R2220 VSS.n1017 VSS.n495 23.5962
R2221 VSS.t197 VSS.n129 23.5962
R2222 VSS.n1261 VSS.n233 23.5962
R2223 VSS.n1299 VSS.n1298 23.4964
R2224 VSS.n1298 VSS.n192 23.4087
R2225 VSS.n1317 VSS.n166 23.3249
R2226 VSS.n1341 VSS.n1340 23.3249
R2227 VSS.n1372 VSS.n100 23.3249
R2228 VSS.n834 VSS.n726 23.3249
R2229 VSS.n867 VSS.n2 23.3249
R2230 VSS.n872 VSS.t2 23.3012
R2231 VSS.t231 VSS.t161 23.3012
R2232 VSS.n1381 VSS.t165 23.3012
R2233 VSS.t86 VSS.t200 23.3012
R2234 VSS.n154 VSS.t153 23.0063
R2235 VSS.n300 VSS.n299 22.8576
R2236 VSS.n299 VSS.n298 22.8576
R2237 VSS.n298 VSS.n297 22.8576
R2238 VSS.n297 VSS.n296 22.8576
R2239 VSS.n296 VSS.n295 22.8576
R2240 VSS.n1226 VSS.n1225 22.8576
R2241 VSS.n1225 VSS.n1224 22.8576
R2242 VSS.n1224 VSS.n1223 22.8576
R2243 VSS.n1223 VSS.n1222 22.8576
R2244 VSS.n514 VSS.n513 22.8576
R2245 VSS.n515 VSS.n514 22.8576
R2246 VSS.n516 VSS.n515 22.8576
R2247 VSS.n517 VSS.n516 22.8576
R2248 VSS.n985 VSS.n517 22.8576
R2249 VSS.n521 VSS.n520 22.8576
R2250 VSS.n520 VSS.n519 22.8576
R2251 VSS.n519 VSS.n518 22.8576
R2252 VSS.n518 VSS.n75 22.8576
R2253 VSS.n473 VSS.n472 22.8576
R2254 VSS.n472 VSS.n471 22.8576
R2255 VSS.n471 VSS.n470 22.8576
R2256 VSS.n470 VSS.n469 22.8576
R2257 VSS.n469 VSS.n468 22.8576
R2258 VSS.n1398 VSS.n1397 22.8576
R2259 VSS.n1397 VSS.n1396 22.8576
R2260 VSS.n1396 VSS.n1395 22.8576
R2261 VSS.n1395 VSS.n1394 22.8576
R2262 VSS.n1037 VSS.n1036 22.8576
R2263 VSS.n1036 VSS.n1035 22.8576
R2264 VSS.n1035 VSS.n1034 22.8576
R2265 VSS.n1034 VSS.n1033 22.8576
R2266 VSS.n1033 VSS.n1032 22.8576
R2267 VSS.n485 VSS.n484 22.8576
R2268 VSS.n486 VSS.n485 22.8576
R2269 VSS.n487 VSS.n486 22.8576
R2270 VSS.n488 VSS.n487 22.8576
R2271 VSS.n1048 VSS.n1047 22.8576
R2272 VSS.n1047 VSS.n1046 22.8576
R2273 VSS.n1046 VSS.n1045 22.8576
R2274 VSS.n1045 VSS.n1044 22.8576
R2275 VSS.n1044 VSS.n1043 22.8576
R2276 VSS.n508 VSS.n456 22.8576
R2277 VSS.n508 VSS.n506 22.8576
R2278 VSS.n506 VSS.n504 22.8576
R2279 VSS.n504 VSS.n502 22.8576
R2280 VSS.n349 VSS.n348 22.8576
R2281 VSS.n350 VSS.n349 22.8576
R2282 VSS.n351 VSS.n350 22.8576
R2283 VSS.n352 VSS.n351 22.8576
R2284 VSS.n1196 VSS.n352 22.8576
R2285 VSS.n1193 VSS.n1192 22.8576
R2286 VSS.n1192 VSS.n1191 22.8576
R2287 VSS.n1191 VSS.n1190 22.8576
R2288 VSS.n1190 VSS.n274 22.8576
R2289 VSS.n292 VSS.n290 22.8576
R2290 VSS.n290 VSS.n288 22.8576
R2291 VSS.n288 VSS.n286 22.8576
R2292 VSS.n286 VSS.n284 22.8576
R2293 VSS.n284 VSS.n223 22.8576
R2294 VSS.n1270 VSS.n1269 22.8576
R2295 VSS.n1269 VSS.n1268 22.8576
R2296 VSS.n1268 VSS.n1267 22.8576
R2297 VSS.n1267 VSS.n209 22.8576
R2298 VSS.n1281 VSS.n1280 22.8576
R2299 VSS.n1280 VSS.n1279 22.8576
R2300 VSS.n1279 VSS.n1278 22.8576
R2301 VSS.n1278 VSS.n1277 22.8576
R2302 VSS.n1277 VSS.n1276 22.8576
R2303 VSS.n1174 VSS.n1173 22.8576
R2304 VSS.n1176 VSS.n1174 22.8576
R2305 VSS.n1176 VSS.n1175 22.8576
R2306 VSS.n1175 VSS.n1166 22.8576
R2307 VSS.n1313 VSS.n170 22.7012
R2308 VSS.n1102 VSS.n411 22.6687
R2309 VSS.t90 VSS.n169 22.4164
R2310 VSS.n164 VSS.n151 22.1254
R2311 VSS.n1351 VSS.n121 22.1254
R2312 VSS.n782 VSS.n98 22.1254
R2313 VSS.n724 VSS.n712 22.1254
R2314 VSS.n335 VSS.n334 22.1254
R2315 VSS.n618 VSS.n604 22.1254
R2316 VSS.t144 VSS.t11 22.1214
R2317 VSS.n807 VSS.n86 22.1214
R2318 VSS.t129 VSS.t108 22.1214
R2319 VSS.n872 VSS.t198 21.8265
R2320 VSS.n1385 VSS.n80 21.8265
R2321 VSS.n1422 VSS.n1421 21.6672
R2322 VSS.n1421 VSS.n29 21.6672
R2323 VSS.n640 VSS.n34 21.6672
R2324 VSS.n34 VSS.n29 21.6672
R2325 VSS.n1136 VSS.n1135 21.6672
R2326 VSS.n1135 VSS.n157 21.6672
R2327 VSS.n1123 VSS.n369 21.6672
R2328 VSS.n369 VSS.n157 21.6672
R2329 VSS.n24 VSS.n9 21.6672
R2330 VSS.n29 VSS.n9 21.6672
R2331 VSS.n924 VSS.n8 21.6672
R2332 VSS.n29 VSS.n8 21.6672
R2333 VSS.n1131 VSS.n1130 21.6672
R2334 VSS.n1131 VSS.n157 21.6672
R2335 VSS.n1079 VSS.n373 21.6672
R2336 VSS.n373 VSS.n157 21.6672
R2337 VSS.n1058 VSS.n439 21.4331
R2338 VSS.n886 VSS.t1 21.2366
R2339 VSS.n1419 VSS.n36 21.2366
R2340 VSS.n1323 VSS.n1322 20.9819
R2341 VSS.n141 VSS.n115 20.9819
R2342 VSS.n1378 VSS.n1377 20.9819
R2343 VSS.n840 VSS.n839 20.9819
R2344 VSS.n341 VSS.n340 20.9819
R2345 VSS.n876 VSS.n611 20.9819
R2346 VSS.n565 VSS.n199 20.7761
R2347 VSS.n1364 VSS.t9 20.6467
R2348 VSS.n430 VSS.t105 20.6467
R2349 VSS.n1302 VSS.n184 20.6467
R2350 VSS.n892 VSS.t148 20.3518
R2351 VSS.n735 VSS.n50 20.3518
R2352 VSS.n1400 VSS.n60 20.1784
R2353 VSS.n789 VSS.t167 20.0568
R2354 VSS.t67 VSS.t72 20.0568
R2355 VSS.t203 VSS.n722 19.7619
R2356 VSS.t53 VSS.n731 19.7619
R2357 VSS.n811 VSS.t172 19.7619
R2358 VSS.n755 VSS.n754 19.6928
R2359 VSS.n756 VSS.n755 19.6928
R2360 VSS.n757 VSS.n756 19.6928
R2361 VSS.n758 VSS.n757 19.6928
R2362 VSS.n759 VSS.n758 19.6928
R2363 VSS.n355 VSS.n354 19.6928
R2364 VSS.n356 VSS.n355 19.6928
R2365 VSS.n357 VSS.n356 19.6928
R2366 VSS.n358 VSS.n357 19.6928
R2367 VSS.n1415 VSS.n1414 19.6928
R2368 VSS.n1414 VSS.n1413 19.6928
R2369 VSS.n1413 VSS.n1412 19.6928
R2370 VSS.n1412 VSS.n1411 19.6928
R2371 VSS.n928 VSS.n926 19.6928
R2372 VSS.n930 VSS.n928 19.6928
R2373 VSS.n932 VSS.n930 19.6928
R2374 VSS.n936 VSS.n932 19.6928
R2375 VSS.n936 VSS.n935 19.6928
R2376 VSS.n15 VSS.n13 19.6928
R2377 VSS.n17 VSS.n15 19.6928
R2378 VSS.n19 VSS.n17 19.6928
R2379 VSS.n21 VSS.n19 19.6928
R2380 VSS.n663 VSS.n662 19.6928
R2381 VSS.n662 VSS.n661 19.6928
R2382 VSS.n661 VSS.n660 19.6928
R2383 VSS.n660 VSS.n659 19.6928
R2384 VSS.n659 VSS.n658 19.6928
R2385 VSS.n656 VSS.n655 19.6928
R2386 VSS.n655 VSS.n654 19.6928
R2387 VSS.n654 VSS.n653 19.6928
R2388 VSS.n653 VSS.n527 19.6928
R2389 VSS.n971 VSS.n970 19.6928
R2390 VSS.n970 VSS.n969 19.6928
R2391 VSS.n969 VSS.n968 19.6928
R2392 VSS.n968 VSS.n967 19.6928
R2393 VSS.n967 VSS.n966 19.6928
R2394 VSS.n963 VSS.n962 19.6928
R2395 VSS.n962 VSS.n961 19.6928
R2396 VSS.n961 VSS.n960 19.6928
R2397 VSS.n960 VSS.n53 19.6928
R2398 VSS.n1244 VSS.n1243 19.6928
R2399 VSS.n1243 VSS.n1242 19.6928
R2400 VSS.n1242 VSS.n1241 19.6928
R2401 VSS.n1241 VSS.n1240 19.6928
R2402 VSS.n1240 VSS.n1239 19.6928
R2403 VSS.n1236 VSS.n1235 19.6928
R2404 VSS.n1235 VSS.n1234 19.6928
R2405 VSS.n1234 VSS.n1233 19.6928
R2406 VSS.n1233 VSS.n179 19.6928
R2407 VSS.n1282 VSS.n211 19.5662
R2408 VSS.n731 VSS.n729 19.4669
R2409 VSS.t10 VSS.t191 19.172
R2410 VSS.t124 VSS.t32 19.172
R2411 VSS.n1213 VSS.n279 19.172
R2412 VSS.n1016 VSS.n1015 18.877
R2413 VSS.n248 VSS.t226 18.877
R2414 VSS.t18 VSS.t103 18.5821
R2415 VSS.n490 VSS.n449 18.4691
R2416 VSS.n1424 VSS.n1423 18.2817
R2417 VSS.n1425 VSS.n1424 18.2817
R2418 VSS.n687 VSS.n28 18.2817
R2419 VSS.n1425 VSS.n28 18.2817
R2420 VSS.n1138 VSS.n1137 18.2817
R2421 VSS.n1138 VSS.n156 18.2817
R2422 VSS.n1141 VSS.n1140 18.2817
R2423 VSS.n1140 VSS.n156 18.2817
R2424 VSS.n1427 VSS.n1426 18.2817
R2425 VSS.n1426 VSS.n1425 18.2817
R2426 VSS.n639 VSS.n27 18.2817
R2427 VSS.n1425 VSS.n27 18.2817
R2428 VSS.n378 VSS.n375 18.2817
R2429 VSS.n378 VSS.n156 18.2817
R2430 VSS.n1125 VSS.n1124 18.2817
R2431 VSS.n1125 VSS.n156 18.2817
R2432 VSS.n765 VSS.t121 17.9922
R2433 VSS.n138 VSS.t55 17.6972
R2434 VSS.n1322 VSS.n159 17.683
R2435 VSS.n1314 VSS.n159 17.683
R2436 VSS.n142 VSS.n141 17.683
R2437 VSS.n1337 VSS.n142 17.683
R2438 VSS.n1377 VSS.n93 17.683
R2439 VSS.n1369 VSS.n93 17.683
R2440 VSS.n839 VSS.n718 17.683
R2441 VSS.n831 VSS.n718 17.683
R2442 VSS.n341 VSS.n238 17.683
R2443 VSS.n242 VSS.n238 17.683
R2444 VSS.n617 VSS.n611 17.683
R2445 VSS.n864 VSS.n617 17.683
R2446 VSS.n522 VSS.n521 17.6005
R2447 VSS.n1042 VSS.n456 17.6005
R2448 VSS.n1194 VSS.n1193 17.6005
R2449 VSS.n1271 VSS.n1270 17.6005
R2450 VSS.n682 VSS.n681 17.4501
R2451 VSS.n1150 VSS.n1149 17.4501
R2452 VSS.n945 VSS.t188 17.4023
R2453 VSS.t243 VSS.n1344 17.4023
R2454 VSS.n1090 VSS.t204 17.4023
R2455 VSS.t109 VSS.t179 17.1074
R2456 VSS.t181 VSS.t188 17.1074
R2457 VSS.t210 VSS.t19 16.8124
R2458 VSS.n764 VSS.n763 16.8124
R2459 VSS.n917 VSS.n538 16.5468
R2460 VSS.n1314 VSS.n1313 16.2314
R2461 VSS.n1337 VSS.n1336 16.2314
R2462 VSS.n1369 VSS.n1368 16.2314
R2463 VSS.n831 VSS.n830 16.2314
R2464 VSS.n864 VSS.n863 16.2314
R2465 VSS.t234 VSS.t117 16.2225
R2466 VSS.t54 VSS.n435 16.2225
R2467 VSS.t153 VSS.t89 16.2225
R2468 VSS.t129 VSS.t3 15.9276
R2469 VSS.t204 VSS.n1067 15.6326
R2470 VSS.n1065 VSS.t194 15.6326
R2471 VSS.n585 VSS.n584 15.6103
R2472 VSS.n588 VSS.n587 15.6103
R2473 VSS.n587 VSS.n577 15.6103
R2474 VSS.n584 VSS.n583 15.6103
R2475 VSS.n921 VSS.n536 15.5157
R2476 VSS.n537 VSS.n536 15.5157
R2477 VSS.n899 VSS.n898 15.5157
R2478 VSS.n899 VSS.n578 15.5157
R2479 VSS.n582 VSS.n572 15.5157
R2480 VSS.n582 VSS.n579 15.5157
R2481 VSS.n589 VSS.n581 15.5157
R2482 VSS.n581 VSS.n580 15.5157
R2483 VSS.n568 VSS.n561 15.5157
R2484 VSS.n567 VSS.n566 15.5157
R2485 VSS.n567 VSS.n559 15.5157
R2486 VSS.n569 VSS.n568 15.5157
R2487 VSS.n912 VSS.n560 15.5157
R2488 VSS.n911 VSS.n910 15.5157
R2489 VSS.n910 VSS.n909 15.5157
R2490 VSS.n571 VSS.n560 15.5157
R2491 VSS.t240 VSS.t52 15.3377
R2492 VSS.n934 VSS.n13 15.1636
R2493 VSS.n657 VSS.n656 15.1636
R2494 VSS.n1171 VSS.n231 15.0862
R2495 VSS.n1001 VSS.n492 15.0862
R2496 VSS.n492 VSS.n491 15.0862
R2497 VSS.n231 VSS.n230 15.0862
R2498 VSS.n1203 VSS.n345 14.9948
R2499 VSS.n1000 VSS.n992 14.9948
R2500 VSS.n1348 VSS.t196 14.7478
R2501 VSS.n1103 VSS.n410 14.7205
R2502 VSS.n918 VSS.n917 14.6737
R2503 VSS.n681 VSS.n441 14.6603
R2504 VSS.n1055 VSS.n441 14.6603
R2505 VSS.n1149 VSS.n201 14.6603
R2506 VSS.n1290 VSS.n201 14.6603
R2507 VSS.t97 VSS.t228 14.4528
R2508 VSS.t101 VSS.t53 14.4528
R2509 VSS.t67 VSS.n118 14.4528
R2510 VSS.t49 VSS.t200 14.4528
R2511 VSS.t121 VSS.t71 14.4528
R2512 VSS.n1246 VSS.n1245 14.2748
R2513 VSS.t82 VSS.t21 14.1579
R2514 VSS.n1103 VSS.n1102 13.7605
R2515 VSS.n1186 VSS.n1169 13.7148
R2516 VSS.n1264 VSS.n229 13.7148
R2517 VSS.n1012 VSS.n459 13.7148
R2518 VSS.n1012 VSS.n497 13.7148
R2519 VSS.n1023 VSS.n489 13.7148
R2520 VSS.n1023 VSS.n1022 13.7148
R2521 VSS.n1186 VSS.n1184 13.7148
R2522 VSS.n1264 VSS.n208 13.7148
R2523 VSS.n1207 VSS.n1206 13.6317
R2524 VSS.n677 VSS.n76 13.6317
R2525 VSS.n995 VSS.n994 13.6317
R2526 VSS.n1170 VSS.n275 13.6317
R2527 VSS.n760 VSS.n354 13.2928
R2528 VSS.n964 VSS.n963 13.2928
R2529 VSS.t239 VSS.t56 13.2731
R2530 VSS.n1437 VSS.n7 13.2731
R2531 VSS.t191 VSS.n36 13.2731
R2532 VSS.n826 VSS.t15 13.2731
R2533 VSS.n1168 VSS.n1167 13.133
R2534 VSS.n501 VSS.n498 13.133
R2535 VSS.n1021 VSS.n1020 13.133
R2536 VSS.n1287 VSS.n1286 13.133
R2537 VSS.n1291 VSS.n1290 13.1163
R2538 VSS.n451 VSS.n450 12.9298
R2539 VSS.n452 VSS.n451 12.9298
R2540 VSS.n453 VSS.n452 12.9298
R2541 VSS.n454 VSS.n453 12.9298
R2542 VSS.n455 VSS.n454 12.9298
R2543 VSS.n1008 VSS.n1007 12.9298
R2544 VSS.n1009 VSS.n1008 12.9298
R2545 VSS.n1010 VSS.n1009 12.9298
R2546 VSS.n1011 VSS.n1010 12.9298
R2547 VSS.n465 VSS.n464 12.9298
R2548 VSS.n466 VSS.n465 12.9298
R2549 VSS.n467 VSS.n466 12.9298
R2550 VSS.n482 VSS.n467 12.9298
R2551 VSS.n1030 VSS.n482 12.9298
R2552 VSS.n1028 VSS.n1027 12.9298
R2553 VSS.n1027 VSS.n1026 12.9298
R2554 VSS.n1026 VSS.n1025 12.9298
R2555 VSS.n1025 VSS.n1024 12.9298
R2556 VSS.n213 VSS.n212 12.9298
R2557 VSS.n214 VSS.n213 12.9298
R2558 VSS.n215 VSS.n214 12.9298
R2559 VSS.n216 VSS.n215 12.9298
R2560 VSS.n217 VSS.n216 12.9298
R2561 VSS.n1179 VSS.n1178 12.9298
R2562 VSS.n1178 VSS.n1177 12.9298
R2563 VSS.n1177 VSS.n1165 12.9298
R2564 VSS.n1187 VSS.n1165 12.9298
R2565 VSS.n306 VSS.n305 12.9298
R2566 VSS.n307 VSS.n306 12.9298
R2567 VSS.n308 VSS.n307 12.9298
R2568 VSS.n309 VSS.n308 12.9298
R2569 VSS.n310 VSS.n309 12.9298
R2570 VSS.n225 VSS.n224 12.9298
R2571 VSS.n226 VSS.n225 12.9298
R2572 VSS.n1266 VSS.n226 12.9298
R2573 VSS.n1266 VSS.n1265 12.9298
R2574 VSS.t2 VSS.n614 12.6832
R2575 VSS.n847 VSS.t225 12.6832
R2576 VSS.n1327 VSS.n151 12.5719
R2577 VSS.n1352 VSS.n1351 12.5719
R2578 VSS.n783 VSS.n782 12.5719
R2579 VSS.n844 VSS.n712 12.5719
R2580 VSS.n336 VSS.n335 12.5719
R2581 VSS.n880 VSS.n604 12.5719
R2582 VSS.t211 VSS.t187 12.0933
R2583 VSS.t187 VSS.t230 12.0933
R2584 VSS.n1063 VSS.n143 12.0661
R2585 VSS.n1361 VSS.n108 12.0661
R2586 VSS.n797 VSS.n796 12.0661
R2587 VSS.n250 VSS.n247 12.0661
R2588 VSS.n855 VSS.n854 12.0661
R2589 VSS.n888 VSS.n597 12.0661
R2590 VSS.n914 VSS.n913 11.9393
R2591 VSS.n915 VSS.n914 11.9393
R2592 VSS.n586 VSS.n541 11.9393
R2593 VSS.n915 VSS.n541 11.9393
R2594 VSS.n917 VSS.n916 11.9393
R2595 VSS.n916 VSS.n915 11.9393
R2596 VSS.n897 VSS.n896 11.9393
R2597 VSS.n896 VSS.n895 11.9393
R2598 VSS.n591 VSS.n590 11.9393
R2599 VSS.n895 VSS.n591 11.9393
R2600 VSS.n894 VSS.n570 11.9393
R2601 VSS.n895 VSS.n894 11.9393
R2602 VSS.n555 VSS.n554 11.9393
R2603 VSS.n556 VSS.n555 11.9393
R2604 VSS.n552 VSS.n551 11.9393
R2605 VSS.n551 VSS.n244 11.9393
R2606 VSS.n651 VSS.n530 11.9393
R2607 VSS.n693 VSS.n530 11.9393
R2608 VSS.n657 VSS.n529 11.9393
R2609 VSS.n625 VSS.n529 11.9393
R2610 VSS.n1420 VSS.n35 11.9393
R2611 VSS.n1420 VSS.n1419 11.9393
R2612 VSS.n651 VSS.n6 11.9393
R2613 VSS.n1437 VSS.n6 11.9393
R2614 VSS.n1403 VSS.n57 11.9393
R2615 VSS.n1403 VSS.n1402 11.9393
R2616 VSS.n965 VSS.n55 11.9393
R2617 VSS.n729 VSS.n55 11.9393
R2618 VSS.n1386 VSS.n79 11.9393
R2619 VSS.n1386 VSS.n1385 11.9393
R2620 VSS.n522 VSS.n77 11.9393
R2621 VSS.n793 VSS.n77 11.9393
R2622 VSS.n1006 VSS.n1005 11.9393
R2623 VSS.n1005 VSS.n495 11.9393
R2624 VSS.n87 VSS.n79 11.9393
R2625 VSS.n1381 VSS.n87 11.9393
R2626 VSS.n1042 VSS.n1041 11.9393
R2627 VSS.n1041 VSS.n96 11.9393
R2628 VSS.n1006 VSS.n458 11.9393
R2629 VSS.n1015 VSS.n458 11.9393
R2630 VSS.n1115 VSS.n394 11.9393
R2631 VSS.n1090 VSS.n394 11.9393
R2632 VSS.n1106 VSS.n393 11.9393
R2633 VSS.n1106 VSS.n1105 11.9393
R2634 VSS.n1134 VSS.n370 11.9393
R2635 VSS.n1134 VSS.n1133 11.9393
R2636 VSS.n1115 VSS.n368 11.9393
R2637 VSS.n1066 VSS.n368 11.9393
R2638 VSS.n1161 VSS.n185 11.9393
R2639 VSS.n1302 VSS.n185 11.9393
R2640 VSS.n762 VSS.n761 11.9393
R2641 VSS.n763 VSS.n762 11.9393
R2642 VSS.n1214 VSS.n278 11.9393
R2643 VSS.n1214 VSS.n1213 11.9393
R2644 VSS.n1194 VSS.n276 11.9393
R2645 VSS.n328 VSS.n276 11.9393
R2646 VSS.n1182 VSS.n1181 11.9393
R2647 VSS.n1182 VSS.n233 11.9393
R2648 VSS.n316 VSS.n278 11.9393
R2649 VSS.n1209 VSS.n316 11.9393
R2650 VSS.n1275 VSS.n1274 11.9393
R2651 VSS.n1274 VSS.n1273 11.9393
R2652 VSS.n1181 VSS.n1180 11.9393
R2653 VSS.n1180 VSS.n235 11.9393
R2654 VSS.n1435 VSS.n11 11.9393
R2655 VSS.n693 VSS.n11 11.9393
R2656 VSS.n934 VSS.n534 11.9393
R2657 VSS.n625 VSS.n534 11.9393
R2658 VSS.n1418 VSS.n1417 11.9393
R2659 VSS.n1419 VSS.n1418 11.9393
R2660 VSS.n1436 VSS.n1435 11.9393
R2661 VSS.n1437 VSS.n1436 11.9393
R2662 VSS.n1401 VSS.n1400 11.9393
R2663 VSS.n1402 VSS.n1401 11.9393
R2664 VSS.n728 VSS.n39 11.9393
R2665 VSS.n729 VSS.n728 11.9393
R2666 VSS.n1384 VSS.n1383 11.9393
R2667 VSS.n1385 VSS.n1384 11.9393
R2668 VSS.n792 VSS.n61 11.9393
R2669 VSS.n793 VSS.n792 11.9393
R2670 VSS.n1029 VSS.n483 11.9393
R2671 VSS.n495 VSS.n483 11.9393
R2672 VSS.n1383 VSS.n1382 11.9393
R2673 VSS.n1382 VSS.n1381 11.9393
R2674 VSS.n1031 VSS.n462 11.9393
R2675 VSS.n462 VSS.n96 11.9393
R2676 VSS.n1029 VSS.n461 11.9393
R2677 VSS.n1015 VSS.n461 11.9393
R2678 VSS.n1089 VSS.n1088 11.9393
R2679 VSS.n1090 VSS.n1089 11.9393
R2680 VSS.n1104 VSS.n1103 11.9393
R2681 VSS.n1105 VSS.n1104 11.9393
R2682 VSS.n1132 VSS.n260 11.9393
R2683 VSS.n1133 VSS.n1132 11.9393
R2684 VSS.n1088 VSS.n374 11.9393
R2685 VSS.n1066 VSS.n374 11.9393
R2686 VSS.n1303 VSS.n183 11.9393
R2687 VSS.n1303 VSS.n1302 11.9393
R2688 VSS.n1238 VSS.n181 11.9393
R2689 VSS.n763 VSS.n181 11.9393
R2690 VSS.n1212 VSS.n1211 11.9393
R2691 VSS.n1213 VSS.n1212 11.9393
R2692 VSS.n327 VSS.n262 11.9393
R2693 VSS.n328 VSS.n327 11.9393
R2694 VSS.n313 VSS.n312 11.9393
R2695 VSS.n313 VSS.n233 11.9393
R2696 VSS.n1211 VSS.n1210 11.9393
R2697 VSS.n1210 VSS.n1209 11.9393
R2698 VSS.n1272 VSS.n1271 11.9393
R2699 VSS.n1273 VSS.n1272 11.9393
R2700 VSS.n312 VSS.n311 11.9393
R2701 VSS.n311 VSS.n235 11.9393
R2702 VSS.n717 VSS.n713 11.9393
R2703 VSS.n714 VSS.n713 11.9393
R2704 VSS.n797 VSS.n788 11.9393
R2705 VSS.n791 VSS.n788 11.9393
R2706 VSS.n805 VSS.n804 11.9393
R2707 VSS.n806 VSS.n805 11.9393
R2708 VSS.n92 VSS.n90 11.9393
R2709 VSS.n1003 VSS.n90 11.9393
R2710 VSS.n431 VSS.n108 11.9393
R2711 VSS.n431 VSS.n430 11.9393
R2712 VSS.n433 VSS.n112 11.9393
R2713 VSS.n434 VSS.n433 11.9393
R2714 VSS.n122 VSS.n117 11.9393
R2715 VSS.n125 VSS.n117 11.9393
R2716 VSS.n145 VSS.n143 11.9393
R2717 VSS.n1062 VSS.n145 11.9393
R2718 VSS.n153 VSS.n149 11.9393
R2719 VSS.n154 VSS.n153 11.9393
R2720 VSS.n158 VSS.n152 11.9393
R2721 VSS.n767 VSS.n152 11.9393
R2722 VSS.n247 VSS.n189 11.9393
R2723 VSS.n189 VSS.n184 11.9393
R2724 VSS.n329 VSS.n193 11.9393
R2725 VSS.n330 VSS.n329 11.9393
R2726 VSS.n339 VSS.n338 11.9393
R2727 VSS.n338 VSS.n279 11.9393
R2728 VSS.n856 VSS.n855 11.9393
R2729 VSS.n857 VSS.n856 11.9393
R2730 VSS.n850 VSS.n849 11.9393
R2731 VSS.n849 VSS.n848 11.9393
R2732 VSS.n875 VSS.n605 11.9393
R2733 VSS.n614 VSS.n605 11.9393
R2734 VSS.n608 VSS.n602 11.9393
R2735 VSS.n608 VSS.n607 11.9393
R2736 VSS.n888 VSS.n887 11.9393
R2737 VSS.n887 VSS.n886 11.9393
R2738 VSS.n1227 VSS.n1226 11.8862
R2739 VSS.n1399 VSS.n1398 11.8862
R2740 VSS VSS.n818 11.7226
R2741 VSS.n779 VSS 11.7226
R2742 VSS.n774 VSS 11.7226
R2743 VSS VSS.n252 11.7226
R2744 VSS.t138 VSS.t223 11.5034
R2745 VSS.t28 VSS.n125 11.5034
R2746 VSS.n720 VSS.n719 11.4711
R2747 VSS.n720 VSS.n36 11.4711
R2748 VSS.n730 VSS.n725 11.4711
R2749 VSS.n731 VSS.n730 11.4711
R2750 VSS.n829 VSS.n727 11.4711
R2751 VSS.n735 VSS.n727 11.4711
R2752 VSS.n781 VSS.n94 11.4711
R2753 VSS.n1016 VSS.n94 11.4711
R2754 VSS.n102 VSS.n99 11.4711
R2755 VSS.n103 VSS.n102 11.4711
R2756 VSS.n1367 VSS.n101 11.4711
R2757 VSS.n811 VSS.n101 11.4711
R2758 VSS.n1350 VSS.n1349 11.4711
R2759 VSS.n1349 VSS.n1348 11.4711
R2760 VSS.n140 VSS.n139 11.4711
R2761 VSS.n139 VSS.n138 11.4711
R2762 VSS.n136 VSS.n132 11.4711
R2763 VSS.n136 VSS.n129 11.4711
R2764 VSS.n161 VSS.n160 11.4711
R2765 VSS.n768 VSS.n161 11.4711
R2766 VSS.n371 VSS.n165 11.4711
R2767 VSS.n372 VSS.n371 11.4711
R2768 VSS.n1312 VSS.n167 11.4711
R2769 VSS.n764 VSS.n167 11.4711
R2770 VSS.n322 VSS.n321 11.4711
R2771 VSS.n321 VSS.n315 11.4711
R2772 VSS.n1259 VSS.n1258 11.4711
R2773 VSS.n1260 VSS.n1259 11.4711
R2774 VSS.n1254 VSS.n243 11.4711
R2775 VSS.n1254 VSS.n1253 11.4711
R2776 VSS.n862 VSS.n620 11.4711
R2777 VSS.n692 VSS.n620 11.4711
R2778 VSS.n870 VSS.n869 11.4711
R2779 VSS.n871 VSS.n870 11.4711
R2780 VSS.n874 VSS.n873 11.4711
R2781 VSS.n873 VSS.n872 11.4711
R2782 VSS.n614 VSS.t95 11.2084
R2783 VSS.n823 VSS.n726 10.9584
R2784 VSS.n810 VSS.n100 10.9584
R2785 VSS.n1341 VSS.n128 10.9584
R2786 VSS.n741 VSS.n166 10.9584
R2787 VSS.n1440 VSS.n2 10.9584
R2788 VSS.n484 VSS.n411 10.7434
R2789 VSS.n622 VSS.n528 10.6369
R2790 VSS.n622 VSS.n531 10.6369
R2791 VSS.n670 VSS.n623 10.6369
R2792 VSS.n623 VSS.n531 10.6369
R2793 VSS.n1092 VSS.n406 10.6369
R2794 VSS.n1093 VSS.n1092 10.6369
R2795 VSS.n1056 VSS.n437 10.6369
R2796 VSS.n1093 VSS.n437 10.6369
R2797 VSS.n947 VSS.n946 10.6369
R2798 VSS.n946 VSS.n945 10.6369
R2799 VSS.n636 VSS.n533 10.6369
R2800 VSS.n945 VSS.n533 10.6369
R2801 VSS.n1108 VSS.n1107 10.6369
R2802 VSS.n1107 VSS.n118 10.6369
R2803 VSS.n407 VSS.n380 10.6369
R2804 VSS.n407 VSS.n118 10.6369
R2805 VSS.n628 VSS.n626 10.6369
R2806 VSS.n626 VSS.n531 10.6369
R2807 VSS.n630 VSS.n627 10.6369
R2808 VSS.n627 VSS.n531 10.6369
R2809 VSS.n1095 VSS.n1094 10.6369
R2810 VSS.n1094 VSS.n1093 10.6369
R2811 VSS.n447 VSS.n436 10.6369
R2812 VSS.n1093 VSS.n436 10.6369
R2813 VSS.n532 VSS.n22 10.6369
R2814 VSS.n945 VSS.n532 10.6369
R2815 VSS.n944 VSS.n943 10.6369
R2816 VSS.n945 VSS.n944 10.6369
R2817 VSS.n421 VSS.n409 10.6369
R2818 VSS.n409 VSS.n118 10.6369
R2819 VSS.n1080 VSS.n408 10.6369
R2820 VSS.n408 VSS.n118 10.6369
R2821 VSS.n848 VSS.n847 10.6185
R2822 VSS.n1402 VSS.t167 10.6185
R2823 VSS.n807 VSS.n806 10.6185
R2824 VSS.n435 VSS.n434 10.6185
R2825 VSS.n155 VSS.n154 10.6185
R2826 VSS.t90 VSS.n168 10.6185
R2827 VSS.n829 VSS.n828 10.3916
R2828 VSS.n1367 VSS.n1366 10.3916
R2829 VSS.n1342 VSS.n132 10.3916
R2830 VSS.n1312 VSS.n1311 10.3916
R2831 VSS.n862 VSS.n861 10.3916
R2832 VSS.t228 VSS.t239 10.3236
R2833 VSS.t203 VSS.t140 10.3236
R2834 VSS.t224 VSS.t171 10.3236
R2835 VSS.n979 VSS.n978 10.2405
R2836 VSS.n980 VSS.n979 10.2405
R2837 VSS.n981 VSS.n980 10.2405
R2838 VSS.n982 VSS.n981 10.2405
R2839 VSS.n983 VSS.n982 10.2405
R2840 VSS.n956 VSS.n955 10.2405
R2841 VSS.n957 VSS.n956 10.2405
R2842 VSS.n959 VSS.n957 10.2405
R2843 VSS.n959 VSS.n958 10.2405
R2844 VSS.n41 VSS.n40 10.2405
R2845 VSS.n42 VSS.n41 10.2405
R2846 VSS.n43 VSS.n42 10.2405
R2847 VSS.n44 VSS.n43 10.2405
R2848 VSS.n255 VSS.n254 10.2405
R2849 VSS.n256 VSS.n255 10.2405
R2850 VSS.n257 VSS.n256 10.2405
R2851 VSS.n258 VSS.n257 10.2405
R2852 VSS.n259 VSS.n258 10.2405
R2853 VSS.n1229 VSS.n1228 10.2405
R2854 VSS.n1230 VSS.n1229 10.2405
R2855 VSS.n1232 VSS.n1230 10.2405
R2856 VSS.n1232 VSS.n1231 10.2405
R2857 VSS.n748 VSS.n747 10.2405
R2858 VSS.n747 VSS.n746 10.2405
R2859 VSS.n746 VSS.n745 10.2405
R2860 VSS.n745 VSS.n744 10.2405
R2861 VSS.n744 VSS.n353 10.2405
R2862 VSS.n1160 VSS.n1159 10.2405
R2863 VSS.n1159 VSS.n1158 10.2405
R2864 VSS.n1158 VSS.n1157 10.2405
R2865 VSS.n1157 VSS.n1156 10.2405
R2866 VSS.t233 VSS.n7 10.0287
R2867 VSS.t139 VSS.t146 10.0287
R2868 VSS.n1007 VSS.n1006 9.95606
R2869 VSS.n1029 VSS.n1028 9.95606
R2870 VSS.n1181 VSS.n1179 9.95606
R2871 VSS.n312 VSS.n224 9.95606
R2872 VSS.n828 VSS.n827 9.91575
R2873 VSS.n827 VSS.n826 9.91575
R2874 VSS.n796 VSS.n795 9.91575
R2875 VSS.n795 VSS.n794 9.91575
R2876 VSS.n1366 VSS.n1365 9.91575
R2877 VSS.n1365 VSS.n1364 9.91575
R2878 VSS.n1362 VSS.n1361 9.91575
R2879 VSS.n1363 VSS.n1362 9.91575
R2880 VSS.n1343 VSS.n1342 9.91575
R2881 VSS.n1344 VSS.n1343 9.91575
R2882 VSS.n1064 VSS.n1063 9.91575
R2883 VSS.n1065 VSS.n1064 9.91575
R2884 VSS.n1311 VSS.n1310 9.91575
R2885 VSS.n1310 VSS.n1309 9.91575
R2886 VSS.n250 VSS.n249 9.91575
R2887 VSS.n249 VSS.n248 9.91575
R2888 VSS.n854 VSS.n696 9.91575
R2889 VSS.n858 VSS.n696 9.91575
R2890 VSS.n861 VSS.n860 9.91575
R2891 VSS.n860 VSS.n7 9.91575
R2892 VSS.n595 VSS.n593 9.91575
R2893 VSS.n593 VSS.t81 9.91575
R2894 VSS.n597 VSS.n594 9.91575
R2895 VSS.n885 VSS.n594 9.91575
R2896 VSS.n562 VSS.n198 9.81228
R2897 VSS.t196 VSS.t28 9.73371
R2898 VSS.n160 VSS.n158 9.65799
R2899 VSS.n1350 VSS.n122 9.65799
R2900 VSS.n781 VSS.n92 9.65799
R2901 VSS.n719 VSS.n717 9.65799
R2902 VSS.n339 VSS.n322 9.65799
R2903 VSS.n875 VSS.n874 9.65799
R2904 VSS.t76 VSS.n825 9.43876
R2905 VSS.t190 VSS.t245 9.14382
R2906 VSS.t220 VSS.t99 9.14382
R2907 VSS.t151 VSS.t88 9.14382
R2908 VSS.n893 VSS.t164 8.84356
R2909 VSS.n1167 VSS 8.81089
R2910 VSS.n501 VSS 8.81089
R2911 VSS.n1020 VSS 8.81089
R2912 VSS.n1286 VSS 8.81089
R2913 VSS.n1275 VSS.n210 8.8005
R2914 VSS.n1173 VSS.n210 8.8005
R2915 VSS.n927 VSS.n925 8.76762
R2916 VSS.n929 VSS.n927 8.76762
R2917 VSS.n931 VSS.n929 8.76762
R2918 VSS.n933 VSS.n931 8.76762
R2919 VSS.n933 VSS.n38 8.76762
R2920 VSS.n14 VSS.n12 8.76762
R2921 VSS.n16 VSS.n14 8.76762
R2922 VSS.n18 VSS.n16 8.76762
R2923 VSS.n20 VSS.n18 8.76762
R2924 VSS.n646 VSS.n645 8.76762
R2925 VSS.n647 VSS.n646 8.76762
R2926 VSS.n648 VSS.n647 8.76762
R2927 VSS.n649 VSS.n648 8.76762
R2928 VSS.n650 VSS.n649 8.76762
R2929 VSS.n954 VSS.n953 8.76762
R2930 VSS.n953 VSS.n952 8.76762
R2931 VSS.n952 VSS.n951 8.76762
R2932 VSS.n951 VSS.n950 8.76762
R2933 VSS.n384 VSS.n382 8.76762
R2934 VSS.n386 VSS.n384 8.76762
R2935 VSS.n388 VSS.n386 8.76762
R2936 VSS.n390 VSS.n388 8.76762
R2937 VSS.n392 VSS.n390 8.76762
R2938 VSS.n398 VSS.n395 8.76762
R2939 VSS.n400 VSS.n398 8.76762
R2940 VSS.n402 VSS.n400 8.76762
R2941 VSS.n404 VSS.n402 8.76762
R2942 VSS.n1077 VSS.n1075 8.76762
R2943 VSS.n1075 VSS.n1073 8.76762
R2944 VSS.n1073 VSS.n1071 8.76762
R2945 VSS.n1071 VSS.n1069 8.76762
R2946 VSS.n1069 VSS.n1068 8.76762
R2947 VSS.n415 VSS.n261 8.76762
R2948 VSS.n416 VSS.n415 8.76762
R2949 VSS.n417 VSS.n416 8.76762
R2950 VSS.n417 VSS.n376 8.76762
R2951 VSS.n1328 VSS.n1327 8.75442
R2952 VSS.n1352 VSS.n120 8.75442
R2953 VSS.n784 VSS.n783 8.75442
R2954 VSS.n336 VSS.n333 8.75442
R2955 VSS.n845 VSS.n844 8.75442
R2956 VSS.n881 VSS.n880 8.75442
R2957 VSS.n898 VSS.n897 8.68898
R2958 VSS.n823 VSS.n822 8.64404
R2959 VSS.n810 VSS.n780 8.64404
R2960 VSS.n775 VSS.n128 8.64404
R2961 VSS.n741 VSS.n740 8.64404
R2962 VSS.n1441 VSS.n1440 8.64404
R2963 VSS.n586 VSS.n585 8.58587
R2964 VSS.t33 VSS.n885 8.55393
R2965 VSS.n607 VSS.t26 8.55393
R2966 VSS.t213 VSS.t231 8.55393
R2967 VSS.n794 VSS.n793 8.55393
R2968 VSS.n1364 VSS.t222 8.55393
R2969 VSS.n590 VSS.n579 8.53383
R2970 VSS.n293 VSS.n291 8.47732
R2971 VSS.n291 VSS.n289 8.47732
R2972 VSS.n289 VSS.n287 8.47732
R2973 VSS.n287 VSS.n285 8.47732
R2974 VSS.n285 VSS.n282 8.47732
R2975 VSS.n264 VSS.n263 8.47732
R2976 VSS.n265 VSS.n264 8.47732
R2977 VSS.n265 VSS.n227 8.47732
R2978 VSS.n228 VSS.n227 8.47732
R2979 VSS.n478 VSS.n477 8.47732
R2980 VSS.n479 VSS.n478 8.47732
R2981 VSS.n480 VSS.n479 8.47732
R2982 VSS.n481 VSS.n480 8.47732
R2983 VSS.n481 VSS.n83 8.47732
R2984 VSS.n63 VSS.n62 8.47732
R2985 VSS.n64 VSS.n63 8.47732
R2986 VSS.n65 VSS.n64 8.47732
R2987 VSS.n66 VSS.n65 8.47732
R2988 VSS.n991 VSS.n990 8.47732
R2989 VSS.n990 VSS.n989 8.47732
R2990 VSS.n989 VSS.n988 8.47732
R2991 VSS.n988 VSS.n987 8.47732
R2992 VSS.n987 VSS.n986 8.47732
R2993 VSS.n510 VSS.n509 8.47732
R2994 VSS.n509 VSS.n507 8.47732
R2995 VSS.n507 VSS.n505 8.47732
R2996 VSS.n505 VSS.n503 8.47732
R2997 VSS.n1202 VSS.n1201 8.47732
R2998 VSS.n1201 VSS.n1200 8.47732
R2999 VSS.n1200 VSS.n1199 8.47732
R3000 VSS.n1199 VSS.n1198 8.47732
R3001 VSS.n1198 VSS.n1197 8.47732
R3002 VSS.n1163 VSS.n1162 8.47732
R3003 VSS.n1164 VSS.n1163 8.47732
R3004 VSS.n1189 VSS.n1164 8.47732
R3005 VSS.n1189 VSS.n1188 8.47732
R3006 VSS.n1020 VSS 8.11479
R3007 VSS.n1167 VSS 8.11479
R3008 VSS.n1416 VSS.n1415 8.07435
R3009 VSS.n1237 VSS.n1236 8.07435
R3010 VSS.t93 VSS.t37 7.96403
R3011 VSS.n955 VSS.n57 7.8853
R3012 VSS.n1161 VSS.n1160 7.8853
R3013 VSS.n501 VSS.n500 7.7784
R3014 VSS.n632 VSS.n631 7.75808
R3015 VSS.n633 VSS.n632 7.75808
R3016 VSS.n634 VSS.n633 7.75808
R3017 VSS.n635 VSS.n634 7.75808
R3018 VSS.n652 VSS.n635 7.75808
R3019 VSS.n524 VSS.n523 7.75808
R3020 VSS.n525 VSS.n524 7.75808
R3021 VSS.n526 VSS.n525 7.75808
R3022 VSS.n949 VSS.n526 7.75808
R3023 VSS.n941 VSS.n940 7.75808
R3024 VSS.n940 VSS.n939 7.75808
R3025 VSS.n939 VSS.n938 7.75808
R3026 VSS.n938 VSS.n937 7.75808
R3027 VSS.n937 VSS.n10 7.75808
R3028 VSS.n1434 VSS.n1433 7.75808
R3029 VSS.n1433 VSS.n1432 7.75808
R3030 VSS.n1432 VSS.n1431 7.75808
R3031 VSS.n1431 VSS.n1430 7.75808
R3032 VSS.n1083 VSS.n1082 7.75808
R3033 VSS.n1084 VSS.n1083 7.75808
R3034 VSS.n1085 VSS.n1084 7.75808
R3035 VSS.n1086 VSS.n1085 7.75808
R3036 VSS.n1087 VSS.n1086 7.75808
R3037 VSS.n413 VSS.n412 7.75808
R3038 VSS.n414 VSS.n413 7.75808
R3039 VSS.n418 VSS.n414 7.75808
R3040 VSS.n419 VSS.n418 7.75808
R3041 VSS.n1121 VSS.n1120 7.75808
R3042 VSS.n1120 VSS.n1119 7.75808
R3043 VSS.n1119 VSS.n1118 7.75808
R3044 VSS.n1118 VSS.n1117 7.75808
R3045 VSS.n1117 VSS.n1116 7.75808
R3046 VSS.n1114 VSS.n1113 7.75808
R3047 VSS.n1113 VSS.n1112 7.75808
R3048 VSS.n1112 VSS.n1111 7.75808
R3049 VSS.n1111 VSS.n1110 7.75808
R3050 VSS.n570 VSS.n569 7.75808
R3051 VSS.n911 VSS.n570 7.75808
R3052 VSS.n913 VSS.n559 7.75808
R3053 VSS.n913 VSS.n912 7.75808
R3054 VSS.n606 VSS.t185 7.66909
R3055 VSS.n1066 VSS.n1065 7.66909
R3056 VSS.n372 VSS.t124 7.66909
R3057 VSS.t52 VSS.t58 7.37414
R3058 VSS.t147 VSS.t162 7.37414
R3059 VSS.n1058 VSS.n1057 7.35731
R3060 VSS.n1286 VSS.n1285 7.18131
R3061 VSS.n1416 VSS.n39 7.08973
R3062 VSS.n1238 VSS.n1237 7.08973
R3063 VSS.n858 VSS.t234 7.0792
R3064 VSS.t69 VSS.t244 7.0792
R3065 VSS.t135 VSS.n175 7.0792
R3066 VSS.n588 VSS.n586 7.02489
R3067 VSS.n590 VSS.n589 6.98232
R3068 VSS.n1031 VSS.n411 6.85764
R3069 VSS.n897 VSS.n537 6.82717
R3070 VSS.n1330 VSS.n1329 6.79974
R3071 VSS.n428 VSS.n427 6.79974
R3072 VSS.n803 VSS.n802 6.79974
R3073 VSS.n326 VSS.n325 6.79974
R3074 VSS.n707 VSS.n706 6.79974
R3075 VSS.n883 VSS.n882 6.79974
R3076 VSS.t96 VSS.t156 6.78425
R3077 VSS.t15 VSS.t75 6.78425
R3078 VSS.t226 VSS.t123 6.78425
R3079 VSS.t73 VSS.n187 6.78425
R3080 VSS.t154 VSS.n330 6.78425
R3081 VSS.n819 VSS 6.60261
R3082 VSS.n736 VSS 6.60261
R3083 VSS VSS.n736 6.60261
R3084 VSS.n738 VSS 6.60261
R3085 VSS VSS.n738 6.60261
R3086 VSS.n739 VSS 6.60261
R3087 VSS.n739 VSS 6.60261
R3088 VSS.n819 VSS 6.60261
R3089 VSS.n1211 VSS.n263 6.52765
R3090 VSS.n1383 VSS.n62 6.52765
R3091 VSS.n510 VSS.n79 6.52765
R3092 VSS.n1162 VSS.n278 6.52765
R3093 VSS.n1003 VSS.n495 6.48931
R3094 VSS.n1344 VSS.t208 6.48931
R3095 VSS.t84 VSS.t159 6.19436
R3096 VSS.n651 VSS.n523 5.97383
R3097 VSS.n1435 VSS.n1434 5.97383
R3098 VSS.n1088 VSS.n412 5.97383
R3099 VSS.n1115 VSS.n1114 5.97383
R3100 VSS.n964 VSS.n954 5.91831
R3101 VSS.n760 VSS.n395 5.91831
R3102 VSS.n1017 VSS.n1016 5.89941
R3103 VSS.t19 VSS.t224 5.89941
R3104 VSS.t130 VSS.n1062 5.89941
R3105 VSS.n1227 VSS.n262 5.71479
R3106 VSS.n1399 VSS.n61 5.71479
R3107 VSS.n1425 VSS.n29 5.60447
R3108 VSS.n1391 VSS.n72 5.60447
R3109 VSS.n1363 VSS.t47 5.60447
R3110 VSS.n1219 VSS.n271 5.60447
R3111 VSS.n1399 VSS.n40 5.3253
R3112 VSS.n1228 VSS.n1227 5.3253
R3113 VSS.n892 VSS.t81 5.30952
R3114 VSS.t106 VSS.t173 5.30952
R3115 VSS.t206 VSS.n156 5.30952
R3116 VSS.n331 VSS.t241 5.30952
R3117 VSS.n295 VSS.n262 5.25764
R3118 VSS.n468 VSS.n61 5.25764
R3119 VSS.n1032 VSS.n1031 5.25764
R3120 VSS.n1043 VSS.n1042 5.25764
R3121 VSS.n1271 VSS.n223 5.25764
R3122 VSS.n1276 VSS.n1275 5.25764
R3123 VSS.n701 VSS.t83 5.18221
R3124 VSS.n602 VSS.t189 5.18221
R3125 VSS.n705 VSS.t212 5.18221
R3126 VSS.n850 VSS.t176 5.18221
R3127 VSS.n1297 VSS.t134 5.18221
R3128 VSS.n193 VSS.t74 5.18221
R3129 VSS.n194 VSS.t207 5.18221
R3130 VSS.n149 VSS.t50 5.18221
R3131 VSS.n1357 VSS.t68 5.18221
R3132 VSS.n112 VSS.t219 5.18221
R3133 VSS.n786 VSS.t166 5.18221
R3134 VSS.n804 VSS.t17 5.18221
R3135 VSS.t229 VSS.t225 5.01458
R3136 VSS.t87 VSS.t45 5.01458
R3137 VSS.n985 VSS.n984 4.91479
R3138 VSS.n1196 VSS.n1195 4.91479
R3139 VSS.n1441 VSS 4.78829
R3140 VSS.n871 VSS.t92 4.71963
R3141 VSS.n768 VSS.t87 4.71963
R3142 VSS.n548 VSS.n547 4.55782
R3143 VSS.n761 VSS.n759 4.52973
R3144 VSS.n935 VSS.n934 4.52973
R3145 VSS.n658 VSS.n657 4.52973
R3146 VSS.n966 VSS.n965 4.52973
R3147 VSS.n1239 VSS.n1238 4.52973
R3148 VSS.t1 VSS.t113 4.42469
R3149 VSS.n825 VSS.n735 4.42469
R3150 VSS.t183 VSS.t54 4.42469
R3151 VSS.n1345 VSS.n129 4.42469
R3152 VSS.n765 VSS.n764 4.42469
R3153 VSS.n1253 VSS.n1252 4.42469
R3154 VSS.n1294 VSS.n1293 4.25121
R3155 VSS.n448 VSS.n446 4.20621
R3156 VSS.n597 VSS.t110 4.17407
R3157 VSS.n1063 VSS.t205 4.17407
R3158 VSS.n1361 VSS.t70 4.17407
R3159 VSS.n796 VSS.t168 4.17407
R3160 VSS.n250 VSS.t136 4.17407
R3161 VSS.n854 VSS.t214 4.17407
R3162 VSS.t93 VSS.t159 4.12974
R3163 VSS VSS.n1442 4.03714
R3164 VSS.n1408 VSS.n50 3.83479
R3165 VSS.n1308 VSS.n175 3.83479
R3166 VSS.n331 VSS.t154 3.83479
R3167 VSS.n1416 VSS.n12 3.59502
R3168 VSS.n1237 VSS.n261 3.59502
R3169 VSS.n714 VSS.t10 3.53985
R3170 VSS.n1319 VSS.n164 3.31902
R3171 VSS.n133 VSS.n121 3.31902
R3172 VSS.n1374 VSS.n98 3.31902
R3173 VSS.n836 VSS.n724 3.31902
R3174 VSS.n334 VSS.n239 3.31902
R3175 VSS.n619 VSS.n618 3.31902
R3176 VSS.n1417 VSS.n1416 3.15666
R3177 VSS.n1237 VSS.n260 3.15666
R3178 VSS.n1006 VSS.n455 2.97424
R3179 VSS.n1030 VSS.n1029 2.97424
R3180 VSS.n1181 VSS.n217 2.97424
R3181 VSS.n312 VSS.n310 2.97424
R3182 VSS.n885 VSS.t22 2.94996
R3183 VSS.t140 VSS.n37 2.94996
R3184 VSS.t78 VSS.t182 2.94996
R3185 VSS.n1052 VSS.n103 2.94996
R3186 VSS.n1345 VSS.t242 2.94996
R3187 VSS.n1293 VSS.n198 2.94342
R3188 VSS.n907 VSS.n906 2.65959
R3189 VSS.n906 VSS.n905 2.65959
R3190 VSS.n904 VSS.n903 2.65959
R3191 VSS.n905 VSS.n904 2.65959
R3192 VSS.n540 VSS.n535 2.65959
R3193 VSS.n905 VSS.n540 2.65959
R3194 VSS.n564 VSS.n557 2.65959
R3195 VSS.n905 VSS.n557 2.65959
R3196 VSS.t227 VSS.t181 2.65501
R3197 VSS.t82 VSS.t36 2.65501
R3198 VSS.t175 VSS.n29 2.65501
R3199 VSS.t48 VSS.t72 2.65501
R3200 VSS.t133 VSS.t155 2.65501
R3201 VSS.n1145 VSS.n279 2.65501
R3202 VSS.n1400 VSS.n1399 2.5605
R3203 VSS.n1227 VSS.n183 2.5605
R3204 VSS.n1283 VSS.n1282 2.37582
R3205 VSS.n643 VSS.n642 2.36762
R3206 VSS.n672 VSS.n671 2.36762
R3207 VSS.n366 VSS.n361 2.36762
R3208 VSS.n1128 VSS.n1127 2.36762
R3209 VSS.n692 VSS.n5 2.36007
R3210 VSS.t201 VSS.n104 2.36007
R3211 VSS.t232 VSS.n811 2.36007
R3212 VSS.n259 VSS.n183 2.3557
R3213 VSS.n984 VSS.n983 2.2021
R3214 VSS.n1195 VSS.n353 2.2021
R3215 VSS.t26 VSS.n606 2.06512
R3216 VSS.n1438 VSS.n5 2.06512
R3217 VSS.t128 VSS.t193 2.06512
R3218 VSS.t106 VSS.t182 2.06512
R3219 VSS.n812 VSS.t232 2.06512
R3220 VSS.t80 VSS.t195 2.06512
R3221 VSS.t155 VSS.t41 2.06512
R3222 VSS.t23 VSS.t163 2.06512
R3223 VSS.n1417 VSS.n38 2.01694
R3224 VSS.n650 VSS.n35 2.01694
R3225 VSS.n392 VSS.n370 2.01694
R3226 VSS.n1068 VSS.n260 2.01694
R3227 VSS.n1211 VSS.n282 1.95017
R3228 VSS.n1383 VSS.n83 1.95017
R3229 VSS.n986 VSS.n79 1.95017
R3230 VSS.n1197 VSS.n278 1.95017
R3231 VSS.n674 VSS.n673 1.92927
R3232 VSS.n976 VSS.n975 1.92927
R3233 VSS.n750 VSS.n749 1.92927
R3234 VSS.n1154 VSS.n1153 1.92927
R3235 VSS.n761 VSS.n760 1.87127
R3236 VSS.n965 VSS.n964 1.87127
R3237 VSS.n1221 VSS.n266 1.81543
R3238 VSS.n1393 VSS.n67 1.81543
R3239 VSS.n1389 VSS.n1388 1.81543
R3240 VSS.n1217 VSS.n1216 1.81543
R3241 VSS.n652 VSS.n651 1.78474
R3242 VSS.n1435 VSS.n10 1.78474
R3243 VSS.n1088 VSS.n1087 1.78474
R3244 VSS.n1116 VSS.n1115 1.78474
R3245 VSS.n667 VSS.n625 1.77017
R3246 VSS.t16 VSS.t192 1.77017
R3247 VSS.n1105 VSS.n104 1.77017
R3248 VSS.n347 VSS.n346 1.73764
R3249 VSS.n1124 VSS.n1123 1.73764
R3250 VSS.n512 VSS.n511 1.73764
R3251 VSS.n640 VSS.n639 1.73764
R3252 VSS.n1330 VSS.n148 1.69426
R3253 VSS.n428 VSS.n109 1.69426
R3254 VSS.n802 VSS.n737 1.69426
R3255 VSS.n325 VSS.n251 1.69426
R3256 VSS.n706 VSS.n700 1.69426
R3257 VSS.n883 VSS.n601 1.69426
R3258 VSS.t20 VSS.t109 1.47523
R3259 VSS.n548 VSS.n545 1.32679
R3260 VSS.n550 VSS.n549 1.22171
R3261 VSS.n753 VSS.n752 1.18907
R3262 VSS.n973 VSS.n972 1.18907
R3263 VSS.n791 VSS.t220 1.18028
R3264 VSS.n703 VSS.n597 1.13213
R3265 VSS.n1063 VSS.n111 1.09859
R3266 VSS.n1361 VSS.n1360 1.09859
R3267 VSS.n796 VSS.n704 1.09859
R3268 VSS.n250 VSS.n197 1.09859
R3269 VSS.n854 VSS.n853 1.09859
R3270 VSS.n1049 VSS.n449 1.09764
R3271 VSS.n1246 VSS.n252 1.07839
R3272 VSS.n547 VSS.t216 1.0711
R3273 VSS.n547 VSS.t238 1.0711
R3274 VSS.n1130 VSS.n375 1.04878
R3275 VSS.n1423 VSS.n1422 1.04878
R3276 VSS.n1427 VSS.n24 1.04878
R3277 VSS.n1137 VSS.n1136 1.04878
R3278 VSS.n360 VSS.n359 0.935332
R3279 VSS.n1410 VSS.n45 0.935332
R3280 VSS.n1406 VSS.n1405 0.935332
R3281 VSS.n1306 VSS.n1305 0.935332
R3282 VSS.n945 VSS.n531 0.885337
R3283 VSS.n1093 VSS.n118 0.885337
R3284 VSS.n1285 VSS 0.881258
R3285 VSS.n1205 VSS.n1204 0.877212
R3286 VSS.n997 VSS.n996 0.877212
R3287 VSS.n676 VSS.n675 0.877212
R3288 VSS.n1148 VSS.n1144 0.877212
R3289 VSS.n822 VSS.n818 0.850685
R3290 VSS.n780 VSS.n779 0.850685
R3291 VSS.n775 VSS.n774 0.850685
R3292 VSS.n740 VSS.n252 0.850685
R3293 VSS.n964 VSS.n35 0.833377
R3294 VSS.n760 VSS.n370 0.833377
R3295 VSS.n491 VSS.n490 0.6405
R3296 VSS.n230 VSS.n211 0.6405
R3297 VSS.n1169 VSS.n1168 0.582318
R3298 VSS.n498 VSS.n459 0.582318
R3299 VSS.n1022 VSS.n1021 0.582318
R3300 VSS.n1287 VSS.n208 0.582318
R3301 VSS.n1329 VSS.n1328 0.435717
R3302 VSS.n427 VSS.n120 0.435717
R3303 VSS.n803 VSS.n784 0.435717
R3304 VSS.n333 VSS.n326 0.435717
R3305 VSS.n845 VSS.n707 0.435717
R3306 VSS.n882 VSS.n881 0.435717
R3307 VSS.n703 VSS.n702 0.420942
R3308 VSS.n852 VSS.n851 0.420942
R3309 VSS.n1296 VSS.n1295 0.420942
R3310 VSS.n196 VSS.n195 0.420942
R3311 VSS.n1359 VSS.n1358 0.420942
R3312 VSS.n787 VSS.n110 0.420942
R3313 VSS.n396 VSS.n393 0.3845
R3314 VSS.n984 VSS.n522 0.343357
R3315 VSS.n1195 VSS.n1194 0.343357
R3316 VSS.n549 VSS 0.336687
R3317 VSS.n500 VSS 0.329665
R3318 VSS.t209 VSS.t76 0.295446
R3319 VSS.t16 VSS.t221 0.295446
R3320 VSS.n806 VSS.n80 0.295446
R3321 VSS.t149 VSS.t119 0.295446
R3322 VSS.t206 VSS.n157 0.295446
R3323 VSS.t127 VSS.t120 0.295446
R3324 VSS.n1146 VSS.n315 0.295446
R3325 VSS.t146 VSS.t122 0.295446
R3326 VSS.n1261 VSS.n1260 0.295446
R3327 VSS.t23 VSS.t115 0.295446
R3328 VSS.n1253 VSS.n220 0.295446
R3329 VSS.n1442 VSS.n1441 0.293735
R3330 VSS.n636 VSS.n630 0.274786
R3331 VSS.n447 VSS.n380 0.274786
R3332 VSS VSS.n198 0.190696
R3333 VSS.n690 VSS.n689 0.175842
R3334 VSS.n637 VSS.n23 0.175842
R3335 VSS.n425 VSS.n381 0.175842
R3336 VSS.n1061 VSS.n1060 0.175842
R3337 VSS.n628 VSS.n22 0.168921
R3338 VSS.n947 VSS.n528 0.168921
R3339 VSS.n1108 VSS.n406 0.168921
R3340 VSS.n1095 VSS.n421 0.168921
R3341 VSS.n984 VSS.n57 0.1541
R3342 VSS.n1195 VSS.n1161 0.1541
R3343 VSS.n1294 VSS 0.127278
R3344 VSS.n853 VSS.n703 0.124481
R3345 VSS.n852 VSS.n704 0.124481
R3346 VSS.n1360 VSS.n110 0.124481
R3347 VSS.n1359 VSS.n111 0.124481
R3348 VSS.n197 VSS.n196 0.124481
R3349 VSS.n549 VSS.n548 0.101297
R3350 VSS.n1295 VSS.n1294 0.0995958
R3351 VSS.n1171 VSS.n345 0.0919286
R3352 VSS.n1001 VSS.n1000 0.0919286
R3353 VSS.n1207 VSS.n229 0.0836169
R3354 VSS.n677 VSS.n497 0.0836169
R3355 VSS.n994 VSS.n489 0.0836169
R3356 VSS.n1184 VSS.n1170 0.0836169
R3357 VSS.n948 VSS.n32 0.0780758
R3358 VSS.n1429 VSS.n1428 0.0780758
R3359 VSS.n424 VSS.n423 0.0780758
R3360 VSS.n1109 VSS.n364 0.0780758
R3361 VSS.n1293 VSS.n1292 0.0344416
R3362 VSS.n853 VSS.n852 0.0340432
R3363 VSS.n704 VSS.n110 0.0340432
R3364 VSS.n1360 VSS.n1359 0.0340432
R3365 VSS.n196 VSS.n111 0.0340432
R3366 VSS.n1295 VSS.n197 0.0340432
R3367 VSS.n195 VSS.n149 0.019754
R3368 VSS.n1358 VSS.n112 0.019754
R3369 VSS.n804 VSS.n787 0.019754
R3370 VSS.n1296 VSS.n193 0.019754
R3371 VSS.n851 VSS.n850 0.019754
R3372 VSS.n702 VSS.n602 0.019754
R3373 VSS.n195 VSS.n194 0.0197205
R3374 VSS.n1358 VSS.n1357 0.0197205
R3375 VSS.n787 VSS.n786 0.0197205
R3376 VSS.n1297 VSS.n1296 0.0197205
R3377 VSS.n851 VSS.n705 0.0197205
R3378 VSS.n702 VSS.n701 0.0197205
R3379 a_1031_764.t5 a_1031_764.n1 553.975
R3380 a_1031_764.n6 a_1031_764.t5 553.975
R3381 a_1031_764.n5 a_1031_764.t6 275.969
R3382 a_1031_764.n3 a_1031_764.t7 275.969
R3383 a_1031_764.n4 a_1031_764.t4 275.877
R3384 a_1031_764.n9 a_1031_764.t1 15.8632
R3385 a_1031_764.n10 a_1031_764.n9 13.5228
R3386 a_1031_764.n9 a_1031_764.n8 5.588
R3387 a_1031_764.n7 a_1031_764.n6 2.79633
R3388 a_1031_764.n8 a_1031_764.n7 2.52001
R3389 a_1031_764.n3 a_1031_764.n0 2.34014
R3390 a_1031_764.n2 a_1031_764.n3 2.3327
R3391 a_1031_764.n2 a_1031_764.n4 2.23523
R3392 a_1031_764.n4 a_1031_764.n0 2.23295
R3393 a_1031_764.n5 a_1031_764.n2 2.04972
R3394 a_1031_764.n0 a_1031_764.n5 2.04764
R3395 a_1031_764.n10 a_1031_764.t3 1.84683
R3396 a_1031_764.t0 a_1031_764.n10 1.84683
R3397 a_1031_764.n8 a_1031_764.t2 1.73283
R3398 a_1031_764.n7 a_1031_764.n1 1.29633
R3399 a_1031_764.n6 a_1031_764.n0 0.585777
R3400 a_1031_764.n2 a_1031_764.n1 0.569287
R3401 VDD.n303 VDD.n21 837900
R3402 VDD.n136 VDD.n131 77656.5
R3403 VDD.n137 VDD.n136 77656.5
R3404 VDD.n138 VDD.n131 77656.5
R3405 VDD.n138 VDD.n137 77656.5
R3406 VDD.n135 VDD.n129 40146.5
R3407 VDD.n135 VDD.n130 40146.5
R3408 VDD.n139 VDD.n129 40146.5
R3409 VDD.n139 VDD.n130 40146.5
R3410 VDD.n356 VDD.n324 6594.31
R3411 VDD.n324 VDD.n322 6594.31
R3412 VDD.n323 VDD.n322 6594.31
R3413 VDD.n356 VDD.n323 6594.31
R3414 VDD.n360 VDD.n13 5352.1
R3415 VDD.n320 VDD.n13 5352.1
R3416 VDD.n320 VDD.n12 5352.1
R3417 VDD.n360 VDD.n12 5352.1
R3418 VDD.n286 VDD.n34 5352.1
R3419 VDD.n286 VDD.n35 5352.1
R3420 VDD.n282 VDD.n35 5352.1
R3421 VDD.n282 VDD.n34 5352.1
R3422 VDD.n253 VDD.n56 5352.1
R3423 VDD.n253 VDD.n57 5352.1
R3424 VDD.n248 VDD.n57 5352.1
R3425 VDD.n248 VDD.n56 5352.1
R3426 VDD.n216 VDD.n77 5352.1
R3427 VDD.n218 VDD.n77 5352.1
R3428 VDD.n218 VDD.n76 5352.1
R3429 VDD.n216 VDD.n76 5352.1
R3430 VDD.n96 VDD.n89 5352.1
R3431 VDD.n97 VDD.n89 5352.1
R3432 VDD.n177 VDD.n97 5352.1
R3433 VDD.n177 VDD.n96 5352.1
R3434 VDD.n153 VDD.n113 5352.1
R3435 VDD.n153 VDD.n114 5352.1
R3436 VDD.n149 VDD.n114 5352.1
R3437 VDD.n149 VDD.n113 5352.1
R3438 VDD.n372 VDD.n5 3990
R3439 VDD.n374 VDD.n5 3990
R3440 VDD.n10 VDD.n9 3990
R3441 VDD.n364 VDD.n10 3990
R3442 VDD.n307 VDD.n19 3990
R3443 VDD.n307 VDD.n20 3990
R3444 VDD.n292 VDD.n31 3990
R3445 VDD.n290 VDD.n31 3990
R3446 VDD.n269 VDD.n47 3990
R3447 VDD.n271 VDD.n47 3990
R3448 VDD.n53 VDD.n52 3990
R3449 VDD.n256 VDD.n53 3990
R3450 VDD.n233 VDD.n66 3990
R3451 VDD.n235 VDD.n66 3990
R3452 VDD.n70 VDD.n68 3990
R3453 VDD.n231 VDD.n68 3990
R3454 VDD.n212 VDD.n84 3990
R3455 VDD.n208 VDD.n84 3990
R3456 VDD.n204 VDD.n88 3990
R3457 VDD.n202 VDD.n88 3990
R3458 VDD.n171 VDD.n98 3990
R3459 VDD.n171 VDD.n170 3990
R3460 VDD.n159 VDD.n111 3990
R3461 VDD.n157 VDD.n111 3990
R3462 VDD.n368 VDD.n6 3219.52
R3463 VDD.n368 VDD.n4 3219.52
R3464 VDD.n301 VDD.n23 3219.52
R3465 VDD.n301 VDD.n24 3219.52
R3466 VDD.n260 VDD.n48 3219.52
R3467 VDD.n260 VDD.n46 3219.52
R3468 VDD.n232 VDD.n67 3219.52
R3469 VDD.n67 VDD.n65 3219.52
R3470 VDD.n197 VDD.n83 3219.52
R3471 VDD.n197 VDD.n85 3219.52
R3472 VDD.n167 VDD.n105 3219.52
R3473 VDD.n167 VDD.n99 3219.52
R3474 VDD.n132 VDD.n121 2532.29
R3475 VDD.n142 VDD.n141 2527.6
R3476 VDD.n134 VDD.n133 2462.92
R3477 VDD.n140 VDD.n128 2458.49
R3478 VDD.n350 VDD.n346 1307.07
R3479 VDD.n350 VDD.n347 1307.07
R3480 VDD.n352 VDD.n346 1307.07
R3481 VDD.n352 VDD.n347 1307.07
R3482 VDD.n9 VDD.n4 770.484
R3483 VDD.n374 VDD.n4 770.484
R3484 VDD.n364 VDD.n6 770.484
R3485 VDD.n372 VDD.n6 770.484
R3486 VDD.n292 VDD.n24 770.484
R3487 VDD.n24 VDD.n20 770.484
R3488 VDD.n290 VDD.n23 770.484
R3489 VDD.n23 VDD.n19 770.484
R3490 VDD.n52 VDD.n46 770.484
R3491 VDD.n271 VDD.n46 770.484
R3492 VDD.n256 VDD.n48 770.484
R3493 VDD.n269 VDD.n48 770.484
R3494 VDD.n70 VDD.n65 770.484
R3495 VDD.n235 VDD.n65 770.484
R3496 VDD.n232 VDD.n231 770.484
R3497 VDD.n233 VDD.n232 770.484
R3498 VDD.n204 VDD.n85 770.484
R3499 VDD.n208 VDD.n85 770.484
R3500 VDD.n202 VDD.n83 770.484
R3501 VDD.n212 VDD.n83 770.484
R3502 VDD.n159 VDD.n99 770.484
R3503 VDD.n170 VDD.n99 770.484
R3504 VDD.n157 VDD.n105 770.484
R3505 VDD.n105 VDD.n98 770.484
R3506 VDD.n343 VDD.n342 755.732
R3507 VDD.n342 VDD.n341 749.907
R3508 VDD.n476 VDD.t194 648.668
R3509 VDD.n515 VDD.t99 648.668
R3510 VDD.n554 VDD.t128 648.668
R3511 VDD.n593 VDD.t153 648.668
R3512 VDD.n1003 VDD.t197 648.668
R3513 VDD.n974 VDD.t180 648.668
R3514 VDD.n945 VDD.t56 648.668
R3515 VDD.n916 VDD.t87 648.668
R3516 VDD.n887 VDD.t224 648.668
R3517 VDD.n858 VDD.t124 648.668
R3518 VDD.n829 VDD.t13 648.668
R3519 VDD.n123 VDD.n122 521.471
R3520 VDD.n125 VDD.n124 506.445
R3521 VDD.n148 VDD.n116 457.914
R3522 VDD.n148 VDD.n110 457.914
R3523 VDD.n449 VDD.t95 372.885
R3524 VDD.n431 VDD.t201 372.885
R3525 VDD.n413 VDD.t46 372.885
R3526 VDD.n395 VDD.t191 372.885
R3527 VDD.n631 VDD.t199 372.885
R3528 VDD.n659 VDD.t101 372.885
R3529 VDD.n687 VDD.t54 372.885
R3530 VDD.n715 VDD.t81 372.885
R3531 VDD.n743 VDD.t110 372.885
R3532 VDD.n771 VDD.t93 372.885
R3533 VDD.n799 VDD.t11 372.885
R3534 VDD.t129 VDD.n346 341.101
R3535 VDD.t115 VDD.n347 341.101
R3536 VDD.n467 VDD.n453 321.882
R3537 VDD.n470 VDD.n451 321.882
R3538 VDD.n447 VDD.n446 321.882
R3539 VDD.n484 VDD.n483 321.882
R3540 VDD.n494 VDD.n493 321.882
R3541 VDD.n506 VDD.n438 321.882
R3542 VDD.n509 VDD.n433 321.882
R3543 VDD.n429 VDD.n428 321.882
R3544 VDD.n523 VDD.n522 321.882
R3545 VDD.n533 VDD.n532 321.882
R3546 VDD.n545 VDD.n420 321.882
R3547 VDD.n548 VDD.n415 321.882
R3548 VDD.n411 VDD.n410 321.882
R3549 VDD.n562 VDD.n561 321.882
R3550 VDD.n572 VDD.n571 321.882
R3551 VDD.n584 VDD.n402 321.882
R3552 VDD.n587 VDD.n397 321.882
R3553 VDD.n393 VDD.n392 321.882
R3554 VDD.n601 VDD.n600 321.882
R3555 VDD.n611 VDD.n610 321.882
R3556 VDD.n624 VDD.n384 321.882
R3557 VDD.n627 VDD.n379 321.882
R3558 VDD.n637 VDD.n636 321.882
R3559 VDD.n650 VDD.n640 321.882
R3560 VDD.n642 VDD.n641 321.882
R3561 VDD.n654 VDD.n643 321.882
R3562 VDD.n657 VDD.n648 321.882
R3563 VDD.n665 VDD.n664 321.882
R3564 VDD.n678 VDD.n668 321.882
R3565 VDD.n670 VDD.n669 321.882
R3566 VDD.n682 VDD.n671 321.882
R3567 VDD.n685 VDD.n676 321.882
R3568 VDD.n693 VDD.n692 321.882
R3569 VDD.n706 VDD.n696 321.882
R3570 VDD.n698 VDD.n697 321.882
R3571 VDD.n710 VDD.n699 321.882
R3572 VDD.n713 VDD.n704 321.882
R3573 VDD.n721 VDD.n720 321.882
R3574 VDD.n734 VDD.n724 321.882
R3575 VDD.n726 VDD.n725 321.882
R3576 VDD.n738 VDD.n727 321.882
R3577 VDD.n741 VDD.n732 321.882
R3578 VDD.n749 VDD.n748 321.882
R3579 VDD.n762 VDD.n752 321.882
R3580 VDD.n754 VDD.n753 321.882
R3581 VDD.n766 VDD.n755 321.882
R3582 VDD.n769 VDD.n760 321.882
R3583 VDD.n777 VDD.n776 321.882
R3584 VDD.n790 VDD.n780 321.882
R3585 VDD.n782 VDD.n781 321.882
R3586 VDD.n794 VDD.n783 321.882
R3587 VDD.n797 VDD.n788 321.882
R3588 VDD.n805 VDD.n804 321.882
R3589 VDD.n810 VDD.n808 321.882
R3590 VDD.n376 VDD.n375 303.579
R3591 VDD.n116 VDD.n115 295.428
R3592 VDD.n214 VDD.n80 295.428
R3593 VDD.n215 VDD.n72 295.428
R3594 VDD.n265 VDD.n264 295.401
R3595 VDD.n263 VDD.n49 294.411
R3596 VDD.n362 VDD.n361 289.565
R3597 VDD.n266 VDD.n265 272.565
R3598 VDD.n273 VDD.n30 272.188
R3599 VDD.n457 VDD.n452 271.068
R3600 VDD.n473 VDD.n434 271.068
R3601 VDD.n512 VDD.n416 271.068
R3602 VDD.n551 VDD.n398 271.068
R3603 VDD.n590 VDD.n380 271.068
R3604 VDD.n649 VDD.n635 271.068
R3605 VDD.n677 VDD.n663 271.068
R3606 VDD.n705 VDD.n691 271.068
R3607 VDD.n733 VDD.n719 271.068
R3608 VDD.n761 VDD.n747 271.068
R3609 VDD.n789 VDD.n775 271.068
R3610 VDD.n809 VDD.n803 271.068
R3611 VDD.n816 VDD.n813 271.068
R3612 VDD.n469 VDD.t211 269.426
R3613 VDD.n462 VDD.t236 255.935
R3614 VDD.n501 VDD.t243 255.935
R3615 VDD.n540 VDD.t239 255.935
R3616 VDD.n579 VDD.t248 255.935
R3617 VDD.n619 VDD.t235 255.935
R3618 VDD.n982 VDD.t234 255.935
R3619 VDD.n953 VDD.t238 255.935
R3620 VDD.n924 VDD.t237 255.935
R3621 VDD.n895 VDD.t245 255.935
R3622 VDD.n866 VDD.t240 255.935
R3623 VDD.n837 VDD.t244 255.935
R3624 VDD VDD.n80 250.803
R3625 VDD.n215 VDD 250.803
R3626 VDD VDD.n49 250.803
R3627 VDD.n361 VDD 250.75
R3628 VDD.n102 VDD.n101 248.601
R3629 VDD.n319 VDD.n14 248.601
R3630 VDD.n239 VDD.n238 248.601
R3631 VDD.n219 VDD.n75 248.601
R3632 VDD.n101 VDD.n87 246.88
R3633 VDD.n161 VDD.n110 246.88
R3634 VDD.n319 VDD.n318 246.88
R3635 VDD.n294 VDD.n30 246.88
R3636 VDD.n241 VDD.n239 246.88
R3637 VDD.n221 VDD.n219 246.88
R3638 VDD.n456 VDD.t212 224.672
R3639 VDD.n441 VDD.t221 224.672
R3640 VDD.n423 VDD.t215 224.672
R3641 VDD.n405 VDD.t155 224.672
R3642 VDD.n387 VDD.t203 224.672
R3643 VDD.n646 VDD.t161 224.672
R3644 VDD.n674 VDD.t209 224.672
R3645 VDD.n702 VDD.t206 224.672
R3646 VDD.n730 VDD.t158 224.672
R3647 VDD.n758 VDD.t218 224.672
R3648 VDD.n786 VDD.t105 224.672
R3649 VDD.n463 VDD.t213 224.492
R3650 VDD.n502 VDD.t222 224.492
R3651 VDD.n541 VDD.t216 224.492
R3652 VDD.n580 VDD.t156 224.492
R3653 VDD.n620 VDD.t204 224.492
R3654 VDD.n981 VDD.t162 224.492
R3655 VDD.n952 VDD.t210 224.492
R3656 VDD.n923 VDD.t207 224.492
R3657 VDD.n894 VDD.t159 224.492
R3658 VDD.n865 VDD.t219 224.492
R3659 VDD.n836 VDD.t106 224.492
R3660 VDD.n812 VDD.t10 217.947
R3661 VDD.n332 VDD.n330 202.397
R3662 VDD.n355 VDD.n339 189.969
R3663 VDD.n471 VDD.n470 185
R3664 VDD.n470 VDD.n469 185
R3665 VDD.n451 VDD.n450 185
R3666 VDD.n467 VDD.n466 185
R3667 VDD.n454 VDD.n453 185
R3668 VDD.n510 VDD.n509 185
R3669 VDD.n509 VDD.n508 185
R3670 VDD.n433 VDD.n432 185
R3671 VDD.n506 VDD.n505 185
R3672 VDD.n439 VDD.n438 185
R3673 VDD.n495 VDD.n494 185
R3674 VDD.n493 VDD.n492 185
R3675 VDD.n483 VDD.n442 185
R3676 VDD.n485 VDD.n484 185
R3677 VDD.n482 VDD.n447 185
R3678 VDD.n446 VDD.n445 185
R3679 VDD.n549 VDD.n548 185
R3680 VDD.n548 VDD.n547 185
R3681 VDD.n415 VDD.n414 185
R3682 VDD.n545 VDD.n544 185
R3683 VDD.n421 VDD.n420 185
R3684 VDD.n534 VDD.n533 185
R3685 VDD.n532 VDD.n531 185
R3686 VDD.n522 VDD.n424 185
R3687 VDD.n524 VDD.n523 185
R3688 VDD.n521 VDD.n429 185
R3689 VDD.n428 VDD.n427 185
R3690 VDD.n588 VDD.n587 185
R3691 VDD.n587 VDD.n586 185
R3692 VDD.n397 VDD.n396 185
R3693 VDD.n584 VDD.n583 185
R3694 VDD.n403 VDD.n402 185
R3695 VDD.n573 VDD.n572 185
R3696 VDD.n571 VDD.n570 185
R3697 VDD.n561 VDD.n406 185
R3698 VDD.n563 VDD.n562 185
R3699 VDD.n560 VDD.n411 185
R3700 VDD.n410 VDD.n409 185
R3701 VDD.n628 VDD.n627 185
R3702 VDD.n627 VDD.n626 185
R3703 VDD.n379 VDD.n378 185
R3704 VDD.n624 VDD.n623 185
R3705 VDD.n385 VDD.n384 185
R3706 VDD.n612 VDD.n611 185
R3707 VDD.n610 VDD.n609 185
R3708 VDD.n600 VDD.n388 185
R3709 VDD.n602 VDD.n601 185
R3710 VDD.n599 VDD.n393 185
R3711 VDD.n392 VDD.n391 185
R3712 VDD.n977 VDD.n657 185
R3713 VDD.n657 VDD.n656 185
R3714 VDD.n978 VDD.n648 185
R3715 VDD.n654 VDD.n644 185
R3716 VDD.n986 VDD.n643 185
R3717 VDD.n987 VDD.n642 185
R3718 VDD.n990 VDD.n641 185
R3719 VDD.n991 VDD.n640 185
R3720 VDD.n650 VDD.n638 185
R3721 VDD.n999 VDD.n637 185
R3722 VDD.n1000 VDD.n636 185
R3723 VDD.n948 VDD.n685 185
R3724 VDD.n685 VDD.n684 185
R3725 VDD.n949 VDD.n676 185
R3726 VDD.n682 VDD.n672 185
R3727 VDD.n957 VDD.n671 185
R3728 VDD.n958 VDD.n670 185
R3729 VDD.n961 VDD.n669 185
R3730 VDD.n962 VDD.n668 185
R3731 VDD.n678 VDD.n666 185
R3732 VDD.n970 VDD.n665 185
R3733 VDD.n971 VDD.n664 185
R3734 VDD.n919 VDD.n713 185
R3735 VDD.n713 VDD.n712 185
R3736 VDD.n920 VDD.n704 185
R3737 VDD.n710 VDD.n700 185
R3738 VDD.n928 VDD.n699 185
R3739 VDD.n929 VDD.n698 185
R3740 VDD.n932 VDD.n697 185
R3741 VDD.n933 VDD.n696 185
R3742 VDD.n706 VDD.n694 185
R3743 VDD.n941 VDD.n693 185
R3744 VDD.n942 VDD.n692 185
R3745 VDD.n890 VDD.n741 185
R3746 VDD.n741 VDD.n740 185
R3747 VDD.n891 VDD.n732 185
R3748 VDD.n738 VDD.n728 185
R3749 VDD.n899 VDD.n727 185
R3750 VDD.n900 VDD.n726 185
R3751 VDD.n903 VDD.n725 185
R3752 VDD.n904 VDD.n724 185
R3753 VDD.n734 VDD.n722 185
R3754 VDD.n912 VDD.n721 185
R3755 VDD.n913 VDD.n720 185
R3756 VDD.n861 VDD.n769 185
R3757 VDD.n769 VDD.n768 185
R3758 VDD.n862 VDD.n760 185
R3759 VDD.n766 VDD.n756 185
R3760 VDD.n870 VDD.n755 185
R3761 VDD.n871 VDD.n754 185
R3762 VDD.n874 VDD.n753 185
R3763 VDD.n875 VDD.n752 185
R3764 VDD.n762 VDD.n750 185
R3765 VDD.n883 VDD.n749 185
R3766 VDD.n884 VDD.n748 185
R3767 VDD.n832 VDD.n797 185
R3768 VDD.n797 VDD.n796 185
R3769 VDD.n833 VDD.n788 185
R3770 VDD.n794 VDD.n784 185
R3771 VDD.n841 VDD.n783 185
R3772 VDD.n842 VDD.n782 185
R3773 VDD.n845 VDD.n781 185
R3774 VDD.n846 VDD.n780 185
R3775 VDD.n790 VDD.n778 185
R3776 VDD.n854 VDD.n777 185
R3777 VDD.n855 VDD.n776 185
R3778 VDD.n817 VDD.n808 185
R3779 VDD.n810 VDD.n806 185
R3780 VDD.n825 VDD.n805 185
R3781 VDD.n826 VDD.n804 185
R3782 VDD.n371 VDD.n2 169.095
R3783 VDD.n274 VDD.n272 161.882
R3784 VDD.n351 VDD.t129 154.345
R3785 VDD.n351 VDD.t115 154.345
R3786 VDD.n444 VDD.n443 153.571
R3787 VDD.n426 VDD.n425 153.571
R3788 VDD.n408 VDD.n407 153.571
R3789 VDD.n390 VDD.n389 153.571
R3790 VDD.n995 VDD.n994 153.571
R3791 VDD.n966 VDD.n965 153.571
R3792 VDD.n937 VDD.n936 153.571
R3793 VDD.n908 VDD.n907 153.571
R3794 VDD.n879 VDD.n878 153.571
R3795 VDD.n850 VDD.n849 153.571
R3796 VDD.n821 VDD.n820 153.571
R3797 VDD.n238 VDD.n236 151.46
R3798 VDD.n207 VDD.n75 151.46
R3799 VDD.n103 VDD.n102 151.46
R3800 VDD.n26 VDD.n14 151.41
R3801 VDD.n508 VDD.t220 118.323
R3802 VDD.n547 VDD.t214 118.323
R3803 VDD.n586 VDD.t154 118.323
R3804 VDD.n626 VDD.t202 118.323
R3805 VDD.n656 VDD.t160 118.323
R3806 VDD.n684 VDD.t208 118.323
R3807 VDD.n712 VDD.t205 118.323
R3808 VDD.n740 VDD.t157 118.323
R3809 VDD.n768 VDD.t217 118.323
R3810 VDD.n796 VDD.t104 118.323
R3811 VDD.n812 VDD.t12 117.838
R3812 VDD.t12 VDD.t0 112.624
R3813 VDD.n370 VDD.n369 112.463
R3814 VDD.n300 VDD.n25 112.463
R3815 VDD.n262 VDD.n261 112.463
R3816 VDD.n227 VDD.n226 112.463
R3817 VDD.n196 VDD.n81 112.463
R3818 VDD.n166 VDD.n106 112.463
R3819 VDD.n123 VDD.t242 105.09
R3820 VDD.n122 VDD.t241 105.09
R3821 VDD.n125 VDD.t246 105.088
R3822 VDD.n124 VDD.t247 105.088
R3823 VDD.n355 VDD.n354 101.487
R3824 VDD.n43 VDD.n42 100.648
R3825 VDD.n318 VDD.n317 99.2798
R3826 VDD.n294 VDD.n293 99.2798
R3827 VDD.n241 VDD.n240 99.2798
R3828 VDD.n221 VDD.n220 99.2798
R3829 VDD.n205 VDD.n87 99.2798
R3830 VDD.n161 VDD.n160 99.2798
R3831 VDD.n375 VDD.n3 90.7299
R3832 VDD.n27 VDD.n26 90.7299
R3833 VDD.n272 VDD.n45 90.7299
R3834 VDD.n236 VDD.n64 90.7299
R3835 VDD.n207 VDD.n206 90.7299
R3836 VDD.n107 VDD.n103 90.7299
R3837 VDD.n317 VDD.n3 90.3534
R3838 VDD.n293 VDD.n27 90.3534
R3839 VDD.n240 VDD.n45 90.3534
R3840 VDD.n220 VDD.n64 90.3534
R3841 VDD.n206 VDD.n205 90.3534
R3842 VDD.n160 VDD.n107 90.3534
R3843 VDD.n468 VDD.n467 86.068
R3844 VDD.n468 VDD.n451 86.068
R3845 VDD.n453 VDD.n452 86.068
R3846 VDD.n447 VDD.n435 86.068
R3847 VDD.n483 VDD.n436 86.068
R3848 VDD.n494 VDD.n437 86.068
R3849 VDD.n507 VDD.n506 86.068
R3850 VDD.n507 VDD.n433 86.068
R3851 VDD.n438 VDD.n437 86.068
R3852 VDD.n493 VDD.n436 86.068
R3853 VDD.n484 VDD.n435 86.068
R3854 VDD.n446 VDD.n434 86.068
R3855 VDD.n429 VDD.n417 86.068
R3856 VDD.n522 VDD.n418 86.068
R3857 VDD.n533 VDD.n419 86.068
R3858 VDD.n546 VDD.n545 86.068
R3859 VDD.n546 VDD.n415 86.068
R3860 VDD.n420 VDD.n419 86.068
R3861 VDD.n532 VDD.n418 86.068
R3862 VDD.n523 VDD.n417 86.068
R3863 VDD.n428 VDD.n416 86.068
R3864 VDD.n411 VDD.n399 86.068
R3865 VDD.n561 VDD.n400 86.068
R3866 VDD.n572 VDD.n401 86.068
R3867 VDD.n585 VDD.n584 86.068
R3868 VDD.n585 VDD.n397 86.068
R3869 VDD.n402 VDD.n401 86.068
R3870 VDD.n571 VDD.n400 86.068
R3871 VDD.n562 VDD.n399 86.068
R3872 VDD.n410 VDD.n398 86.068
R3873 VDD.n393 VDD.n381 86.068
R3874 VDD.n600 VDD.n382 86.068
R3875 VDD.n611 VDD.n383 86.068
R3876 VDD.n625 VDD.n624 86.068
R3877 VDD.n625 VDD.n379 86.068
R3878 VDD.n384 VDD.n383 86.068
R3879 VDD.n610 VDD.n382 86.068
R3880 VDD.n601 VDD.n381 86.068
R3881 VDD.n392 VDD.n380 86.068
R3882 VDD.n651 VDD.n637 86.068
R3883 VDD.n652 VDD.n640 86.068
R3884 VDD.n653 VDD.n642 86.068
R3885 VDD.n655 VDD.n654 86.068
R3886 VDD.n655 VDD.n648 86.068
R3887 VDD.n653 VDD.n643 86.068
R3888 VDD.n652 VDD.n641 86.068
R3889 VDD.n651 VDD.n650 86.068
R3890 VDD.n649 VDD.n636 86.068
R3891 VDD.n679 VDD.n665 86.068
R3892 VDD.n680 VDD.n668 86.068
R3893 VDD.n681 VDD.n670 86.068
R3894 VDD.n683 VDD.n682 86.068
R3895 VDD.n683 VDD.n676 86.068
R3896 VDD.n681 VDD.n671 86.068
R3897 VDD.n680 VDD.n669 86.068
R3898 VDD.n679 VDD.n678 86.068
R3899 VDD.n677 VDD.n664 86.068
R3900 VDD.n707 VDD.n693 86.068
R3901 VDD.n708 VDD.n696 86.068
R3902 VDD.n709 VDD.n698 86.068
R3903 VDD.n711 VDD.n710 86.068
R3904 VDD.n711 VDD.n704 86.068
R3905 VDD.n709 VDD.n699 86.068
R3906 VDD.n708 VDD.n697 86.068
R3907 VDD.n707 VDD.n706 86.068
R3908 VDD.n705 VDD.n692 86.068
R3909 VDD.n735 VDD.n721 86.068
R3910 VDD.n736 VDD.n724 86.068
R3911 VDD.n737 VDD.n726 86.068
R3912 VDD.n739 VDD.n738 86.068
R3913 VDD.n739 VDD.n732 86.068
R3914 VDD.n737 VDD.n727 86.068
R3915 VDD.n736 VDD.n725 86.068
R3916 VDD.n735 VDD.n734 86.068
R3917 VDD.n733 VDD.n720 86.068
R3918 VDD.n763 VDD.n749 86.068
R3919 VDD.n764 VDD.n752 86.068
R3920 VDD.n765 VDD.n754 86.068
R3921 VDD.n767 VDD.n766 86.068
R3922 VDD.n767 VDD.n760 86.068
R3923 VDD.n765 VDD.n755 86.068
R3924 VDD.n764 VDD.n753 86.068
R3925 VDD.n763 VDD.n762 86.068
R3926 VDD.n761 VDD.n748 86.068
R3927 VDD.n791 VDD.n777 86.068
R3928 VDD.n792 VDD.n780 86.068
R3929 VDD.n793 VDD.n782 86.068
R3930 VDD.n795 VDD.n794 86.068
R3931 VDD.n795 VDD.n788 86.068
R3932 VDD.n793 VDD.n783 86.068
R3933 VDD.n792 VDD.n781 86.068
R3934 VDD.n791 VDD.n790 86.068
R3935 VDD.n789 VDD.n776 86.068
R3936 VDD.n811 VDD.n805 86.068
R3937 VDD.n813 VDD.n808 86.068
R3938 VDD.n811 VDD.n810 86.068
R3939 VDD.n809 VDD.n804 86.068
R3940 VDD.n508 VDD.t193 77.2863
R3941 VDD.n547 VDD.t98 77.2863
R3942 VDD.n586 VDD.t127 77.2863
R3943 VDD.n626 VDD.t152 77.2863
R3944 VDD.n656 VDD.t196 77.2863
R3945 VDD.n684 VDD.t179 77.2863
R3946 VDD.n712 VDD.t55 77.2863
R3947 VDD.n740 VDD.t86 77.2863
R3948 VDD.n768 VDD.t223 77.2863
R3949 VDD.n796 VDD.t123 77.2863
R3950 VDD.n344 VDD.n343 74.3011
R3951 VDD.t193 VDD.t107 73.8666
R3952 VDD.t98 VDD.t96 73.8666
R3953 VDD.t127 VDD.t31 73.8666
R3954 VDD.t152 VDD.t41 73.8666
R3955 VDD.t196 VDD.t102 73.8666
R3956 VDD.t179 VDD.t113 73.8666
R3957 VDD.t55 VDD.t8 73.8666
R3958 VDD.t86 VDD.t88 73.8666
R3959 VDD.t223 VDD.t188 73.8666
R3960 VDD.t123 VDD.t84 73.8666
R3961 VDD.n323 VDD.t137 73.412
R3962 VDD.t35 VDD.n324 73.412
R3963 VDD.n341 VDD.n339 70.8706
R3964 VDD.n267 VDD.n266 69.8346
R3965 VDD.n8 VDD.n3 68.9008
R3966 VDD.n299 VDD.n27 68.9008
R3967 VDD.n51 VDD.n45 68.9008
R3968 VDD.n225 VDD.n64 68.9008
R3969 VDD.n206 VDD.n86 68.9008
R3970 VDD.n165 VDD.n107 68.9008
R3971 VDD.t137 VDD.t184 68.2355
R3972 VDD.t184 VDD.t186 68.2355
R3973 VDD.t186 VDD.t76 68.2355
R3974 VDD.t76 VDD.t78 68.2355
R3975 VDD.t78 VDD.t37 68.2355
R3976 VDD.t74 VDD.t39 68.2355
R3977 VDD.t131 VDD.t74 68.2355
R3978 VDD.t139 VDD.t131 68.2355
R3979 VDD.t141 VDD.t139 68.2355
R3980 VDD.t171 VDD.n5 60.7854
R3981 VDD.t82 VDD.n149 59.9455
R3982 VDD.n152 VDD.t62 56.8621
R3983 VDD.n151 VDD.t43 56.8621
R3984 VDD.t6 VDD.n168 56.8621
R3985 VDD.n172 VDD.t4 56.8621
R3986 VDD.n176 VDD.t169 56.8621
R3987 VDD.t177 VDD.n174 56.8621
R3988 VDD.n173 VDD.t135 56.8621
R3989 VDD.n198 VDD.t58 56.8621
R3990 VDD.t133 VDD.n210 56.8621
R3991 VDD.n209 VDD.t117 56.8621
R3992 VDD.t119 VDD.n79 56.8621
R3993 VDD.n78 VDD.t15 56.8621
R3994 VDD.n71 VDD.t111 56.8621
R3995 VDD.t29 VDD.n58 56.8621
R3996 VDD.t143 VDD.n249 56.8621
R3997 VDD.n252 VDD.t145 56.8621
R3998 VDD.n251 VDD.t60 56.8621
R3999 VDD.n259 VDD.t47 56.8621
R4000 VDD.t49 VDD.n36 56.8621
R4001 VDD.t70 VDD.n283 56.8621
R4002 VDD.n285 VDD.t21 56.8621
R4003 VDD.t23 VDD.n32 56.8492
R4004 VDD.n306 VDD.t90 56.8492
R4005 VDD.n305 VDD.t226 56.8492
R4006 VDD.t230 VDD.n358 56.8492
R4007 VDD.n321 VDD.t163 56.8492
R4008 VDD.n367 VDD.t173 56.8492
R4009 VDD.t2 VDD.n104 56.2135
R4010 VDD.n199 VDD.t51 56.2135
R4011 VDD.t66 VDD.n229 56.2135
R4012 VDD.n258 VDD.t182 56.2135
R4013 VDD.t121 VDD.n22 56.2007
R4014 VDD.n366 VDD.t17 56.2007
R4015 VDD.t33 VDD.t82 55.7811
R4016 VDD.t62 VDD.t64 55.7811
R4017 VDD.t169 VDD.t167 55.7811
R4018 VDD.t175 VDD.t177 55.7811
R4019 VDD.t117 VDD.t149 55.7811
R4020 VDD.t147 VDD.t119 55.7811
R4021 VDD.t25 VDD.t143 55.7811
R4022 VDD.t145 VDD.t27 55.7811
R4023 VDD.t72 VDD.t70 55.7811
R4024 VDD.t21 VDD.t19 55.7811
R4025 VDD.t226 VDD.t232 55.7684
R4026 VDD.t228 VDD.t230 55.7684
R4027 VDD.n349 VDD.n348 53.5863
R4028 VDD.n345 VDD.n344 53.3212
R4029 VDD.n349 VDD.n340 51.3524
R4030 VDD.n362 VDD 50.4861
R4031 VDD.t68 VDD.n303 50.3646
R4032 VDD.n469 VDD.n468 49.4675
R4033 VDD.n469 VDD.n452 49.4675
R4034 VDD.n508 VDD.n507 49.4675
R4035 VDD.n508 VDD.n437 49.4675
R4036 VDD.n508 VDD.n436 49.4675
R4037 VDD.n508 VDD.n435 49.4675
R4038 VDD.n508 VDD.n434 49.4675
R4039 VDD.n547 VDD.n546 49.4675
R4040 VDD.n547 VDD.n419 49.4675
R4041 VDD.n547 VDD.n418 49.4675
R4042 VDD.n547 VDD.n417 49.4675
R4043 VDD.n547 VDD.n416 49.4675
R4044 VDD.n586 VDD.n585 49.4675
R4045 VDD.n586 VDD.n401 49.4675
R4046 VDD.n586 VDD.n400 49.4675
R4047 VDD.n586 VDD.n399 49.4675
R4048 VDD.n586 VDD.n398 49.4675
R4049 VDD.n626 VDD.n625 49.4675
R4050 VDD.n626 VDD.n383 49.4675
R4051 VDD.n626 VDD.n382 49.4675
R4052 VDD.n626 VDD.n381 49.4675
R4053 VDD.n626 VDD.n380 49.4675
R4054 VDD.n656 VDD.n655 49.4675
R4055 VDD.n656 VDD.n653 49.4675
R4056 VDD.n656 VDD.n652 49.4675
R4057 VDD.n656 VDD.n651 49.4675
R4058 VDD.n656 VDD.n649 49.4675
R4059 VDD.n684 VDD.n683 49.4675
R4060 VDD.n684 VDD.n681 49.4675
R4061 VDD.n684 VDD.n680 49.4675
R4062 VDD.n684 VDD.n679 49.4675
R4063 VDD.n684 VDD.n677 49.4675
R4064 VDD.n712 VDD.n711 49.4675
R4065 VDD.n712 VDD.n709 49.4675
R4066 VDD.n712 VDD.n708 49.4675
R4067 VDD.n712 VDD.n707 49.4675
R4068 VDD.n712 VDD.n705 49.4675
R4069 VDD.n740 VDD.n739 49.4675
R4070 VDD.n740 VDD.n737 49.4675
R4071 VDD.n740 VDD.n736 49.4675
R4072 VDD.n740 VDD.n735 49.4675
R4073 VDD.n740 VDD.n733 49.4675
R4074 VDD.n768 VDD.n767 49.4675
R4075 VDD.n768 VDD.n765 49.4675
R4076 VDD.n768 VDD.n764 49.4675
R4077 VDD.n768 VDD.n763 49.4675
R4078 VDD.n768 VDD.n761 49.4675
R4079 VDD.n796 VDD.n795 49.4675
R4080 VDD.n796 VDD.n793 49.4675
R4081 VDD.n796 VDD.n792 49.4675
R4082 VDD.n796 VDD.n791 49.4675
R4083 VDD.n796 VDD.n789 49.4675
R4084 VDD.n813 VDD.n812 49.4675
R4085 VDD.n812 VDD.n811 49.4675
R4086 VDD.n812 VDD.n809 49.4675
R4087 VDD.n363 VDD.n11 46.2601
R4088 VDD.n289 VDD.n287 46.2601
R4089 VDD.n255 VDD.n254 46.2601
R4090 VDD.n181 VDD.n69 46.2601
R4091 VDD.n201 VDD.n195 46.2601
R4092 VDD.n156 VDD.n154 46.2601
R4093 VDD VDD.n263 45.8771
R4094 VDD.n115 VDD 44.8603
R4095 VDD VDD.n214 44.8603
R4096 VDD.n72 VDD 44.8603
R4097 VDD.n264 VDD 44.6517
R4098 VDD.n318 VDD.n316 43.4356
R4099 VDD.n295 VDD.n294 43.4356
R4100 VDD.n242 VDD.n241 43.4356
R4101 VDD.n222 VDD.n221 43.4356
R4102 VDD.n191 VDD.n87 43.4356
R4103 VDD.n162 VDD.n161 43.4356
R4104 VDD.n176 VDD.n172 42.3765
R4105 VDD.n210 VDD.n209 42.3765
R4106 VDD.n249 VDD.n58 42.3765
R4107 VDD.n283 VDD.n36 42.3765
R4108 VDD.n306 VDD.n305 42.3668
R4109 VDD.n275 VDD.n274 40.973
R4110 VDD.n309 VDD.n17 40.8986
R4111 VDD.n247 VDD.n59 40.8986
R4112 VDD.n213 VDD.n82 40.8986
R4113 VDD.n178 VDD.n94 40.8986
R4114 VDD.n277 VDD.n276 40.689
R4115 VDD.n18 VDD.n14 39.3388
R4116 VDD.n238 VDD.n237 39.3388
R4117 VDD.n188 VDD.n75 39.3388
R4118 VDD.n102 VDD.n100 39.3388
R4119 VDD.n457 VDD.n454 36.1417
R4120 VDD.n466 VDD.n454 36.1417
R4121 VDD.n466 VDD.n450 36.1417
R4122 VDD.n471 VDD.n450 36.1417
R4123 VDD.n473 VDD.n445 36.1417
R4124 VDD.n482 VDD.n445 36.1417
R4125 VDD.n485 VDD.n482 36.1417
R4126 VDD.n485 VDD.n442 36.1417
R4127 VDD.n492 VDD.n442 36.1417
R4128 VDD.n495 VDD.n439 36.1417
R4129 VDD.n505 VDD.n439 36.1417
R4130 VDD.n505 VDD.n432 36.1417
R4131 VDD.n510 VDD.n432 36.1417
R4132 VDD.n512 VDD.n427 36.1417
R4133 VDD.n521 VDD.n427 36.1417
R4134 VDD.n524 VDD.n521 36.1417
R4135 VDD.n524 VDD.n424 36.1417
R4136 VDD.n531 VDD.n424 36.1417
R4137 VDD.n534 VDD.n421 36.1417
R4138 VDD.n544 VDD.n421 36.1417
R4139 VDD.n544 VDD.n414 36.1417
R4140 VDD.n549 VDD.n414 36.1417
R4141 VDD.n551 VDD.n409 36.1417
R4142 VDD.n560 VDD.n409 36.1417
R4143 VDD.n563 VDD.n560 36.1417
R4144 VDD.n563 VDD.n406 36.1417
R4145 VDD.n570 VDD.n406 36.1417
R4146 VDD.n573 VDD.n403 36.1417
R4147 VDD.n583 VDD.n403 36.1417
R4148 VDD.n583 VDD.n396 36.1417
R4149 VDD.n588 VDD.n396 36.1417
R4150 VDD.n590 VDD.n391 36.1417
R4151 VDD.n599 VDD.n391 36.1417
R4152 VDD.n602 VDD.n599 36.1417
R4153 VDD.n602 VDD.n388 36.1417
R4154 VDD.n609 VDD.n388 36.1417
R4155 VDD.n612 VDD.n385 36.1417
R4156 VDD.n623 VDD.n385 36.1417
R4157 VDD.n623 VDD.n378 36.1417
R4158 VDD.n628 VDD.n378 36.1417
R4159 VDD.n1000 VDD.n635 36.1417
R4160 VDD.n1000 VDD.n999 36.1417
R4161 VDD.n999 VDD.n638 36.1417
R4162 VDD.n991 VDD.n638 36.1417
R4163 VDD.n991 VDD.n990 36.1417
R4164 VDD.n987 VDD.n986 36.1417
R4165 VDD.n986 VDD.n644 36.1417
R4166 VDD.n978 VDD.n644 36.1417
R4167 VDD.n978 VDD.n977 36.1417
R4168 VDD.n971 VDD.n663 36.1417
R4169 VDD.n971 VDD.n970 36.1417
R4170 VDD.n970 VDD.n666 36.1417
R4171 VDD.n962 VDD.n666 36.1417
R4172 VDD.n962 VDD.n961 36.1417
R4173 VDD.n958 VDD.n957 36.1417
R4174 VDD.n957 VDD.n672 36.1417
R4175 VDD.n949 VDD.n672 36.1417
R4176 VDD.n949 VDD.n948 36.1417
R4177 VDD.n942 VDD.n691 36.1417
R4178 VDD.n942 VDD.n941 36.1417
R4179 VDD.n941 VDD.n694 36.1417
R4180 VDD.n933 VDD.n694 36.1417
R4181 VDD.n933 VDD.n932 36.1417
R4182 VDD.n929 VDD.n928 36.1417
R4183 VDD.n928 VDD.n700 36.1417
R4184 VDD.n920 VDD.n700 36.1417
R4185 VDD.n920 VDD.n919 36.1417
R4186 VDD.n913 VDD.n719 36.1417
R4187 VDD.n913 VDD.n912 36.1417
R4188 VDD.n912 VDD.n722 36.1417
R4189 VDD.n904 VDD.n722 36.1417
R4190 VDD.n904 VDD.n903 36.1417
R4191 VDD.n900 VDD.n899 36.1417
R4192 VDD.n899 VDD.n728 36.1417
R4193 VDD.n891 VDD.n728 36.1417
R4194 VDD.n891 VDD.n890 36.1417
R4195 VDD.n884 VDD.n747 36.1417
R4196 VDD.n884 VDD.n883 36.1417
R4197 VDD.n883 VDD.n750 36.1417
R4198 VDD.n875 VDD.n750 36.1417
R4199 VDD.n875 VDD.n874 36.1417
R4200 VDD.n871 VDD.n870 36.1417
R4201 VDD.n870 VDD.n756 36.1417
R4202 VDD.n862 VDD.n756 36.1417
R4203 VDD.n862 VDD.n861 36.1417
R4204 VDD.n855 VDD.n775 36.1417
R4205 VDD.n855 VDD.n854 36.1417
R4206 VDD.n854 VDD.n778 36.1417
R4207 VDD.n846 VDD.n778 36.1417
R4208 VDD.n846 VDD.n845 36.1417
R4209 VDD.n842 VDD.n841 36.1417
R4210 VDD.n841 VDD.n784 36.1417
R4211 VDD.n833 VDD.n784 36.1417
R4212 VDD.n833 VDD.n832 36.1417
R4213 VDD.n826 VDD.n803 36.1417
R4214 VDD.n826 VDD.n825 36.1417
R4215 VDD.n825 VDD.n806 36.1417
R4216 VDD.n817 VDD.n806 36.1417
R4217 VDD.n817 VDD.n816 36.1417
R4218 VDD.n357 VDD.t37 34.118
R4219 VDD.n357 VDD.t39 34.118
R4220 VDD.n351 VDD.t141 34.118
R4221 VDD.n351 VDD.t35 34.118
R4222 VDD.n267 VDD.n37 32.5786
R4223 VDD.n150 VDD.t33 27.8908
R4224 VDD.t64 VDD.n150 27.8908
R4225 VDD.n158 VDD.t43 27.8908
R4226 VDD.n158 VDD.t2 27.8908
R4227 VDD.n169 VDD.t6 27.8908
R4228 VDD.n169 VDD.t4 27.8908
R4229 VDD.t167 VDD.n175 27.8908
R4230 VDD.n175 VDD.t175 27.8908
R4231 VDD.n203 VDD.t135 27.8908
R4232 VDD.n203 VDD.t51 27.8908
R4233 VDD.n211 VDD.t58 27.8908
R4234 VDD.n211 VDD.t133 27.8908
R4235 VDD.n217 VDD.t149 27.8908
R4236 VDD.n217 VDD.t147 27.8908
R4237 VDD.n230 VDD.t15 27.8908
R4238 VDD.n230 VDD.t66 27.8908
R4239 VDD.n234 VDD.t111 27.8908
R4240 VDD.n234 VDD.t29 27.8908
R4241 VDD.n250 VDD.t25 27.8908
R4242 VDD.t27 VDD.n250 27.8908
R4243 VDD.n257 VDD.t60 27.8908
R4244 VDD.t182 VDD.n257 27.8908
R4245 VDD.n270 VDD.t47 27.8908
R4246 VDD.n270 VDD.t49 27.8908
R4247 VDD.n284 VDD.t72 27.8908
R4248 VDD.t19 VDD.n284 27.8908
R4249 VDD.n291 VDD.t23 27.8845
R4250 VDD.n291 VDD.t121 27.8845
R4251 VDD.n304 VDD.t68 27.8845
R4252 VDD.t90 VDD.n304 27.8845
R4253 VDD.n359 VDD.t232 27.8845
R4254 VDD.n359 VDD.t228 27.8845
R4255 VDD.n365 VDD.t163 27.8845
R4256 VDD.t17 VDD.n365 27.8845
R4257 VDD.n373 VDD.t173 27.8845
R4258 VDD.n373 VDD.t171 27.8845
R4259 VDD.n330 VDD.t130 27.6955
R4260 VDD.n330 VDD.t116 27.6955
R4261 VDD.n354 VDD.n353 26.8576
R4262 VDD.n348 VDD.n347 26.4291
R4263 VDD.n346 VDD.n340 26.4291
R4264 VDD.n353 VDD.n345 26.2862
R4265 VDD.n152 VDD.n151 25.945
R4266 VDD.n174 VDD.n173 25.945
R4267 VDD.n79 VDD.n78 25.945
R4268 VDD.n252 VDD.n251 25.945
R4269 VDD.n143 VDD.n120 24.6841
R4270 VDD.t220 VDD.t94 24.6225
R4271 VDD.t214 VDD.t200 24.6225
R4272 VDD.t154 VDD.t45 24.6225
R4273 VDD.t202 VDD.t190 24.6225
R4274 VDD.t160 VDD.t198 24.6225
R4275 VDD.t208 VDD.t100 24.6225
R4276 VDD.t205 VDD.t53 24.6225
R4277 VDD.t157 VDD.t80 24.6225
R4278 VDD.t217 VDD.t109 24.6225
R4279 VDD.t104 VDD.t92 24.6225
R4280 VDD.n127 VDD.n119 24.2261
R4281 VDD.n443 VDD.t192 23.5572
R4282 VDD.n425 VDD.t97 23.5572
R4283 VDD.n407 VDD.t126 23.5572
R4284 VDD.n389 VDD.t151 23.5572
R4285 VDD.n994 VDD.t195 23.5572
R4286 VDD.n965 VDD.t181 23.5572
R4287 VDD.n936 VDD.t57 23.5572
R4288 VDD.n907 VDD.t89 23.5572
R4289 VDD.n878 VDD.t225 23.5572
R4290 VDD.n849 VDD.t125 23.5572
R4291 VDD.n820 VDD.t14 23.5572
R4292 VDD.n357 VDD.n321 23.3452
R4293 VDD.n144 VDD.n119 22.9279
R4294 VDD.n348 VDD.n345 21.5863
R4295 VDD.n276 VDD.n275 20.8005
R4296 VDD.n98 VDD.n94 20.5561
R4297 VDD.n169 VDD.n98 20.5561
R4298 VDD.n157 VDD.n156 20.5561
R4299 VDD.n158 VDD.n157 20.5561
R4300 VDD.n170 VDD.n103 20.5561
R4301 VDD.n170 VDD.n169 20.5561
R4302 VDD.n160 VDD.n159 20.5561
R4303 VDD.n159 VDD.n158 20.5561
R4304 VDD.n213 VDD.n212 20.5561
R4305 VDD.n212 VDD.n211 20.5561
R4306 VDD.n202 VDD.n201 20.5561
R4307 VDD.n203 VDD.n202 20.5561
R4308 VDD.n208 VDD.n207 20.5561
R4309 VDD.n211 VDD.n208 20.5561
R4310 VDD.n205 VDD.n204 20.5561
R4311 VDD.n204 VDD.n203 20.5561
R4312 VDD.n233 VDD.n59 20.5561
R4313 VDD.n234 VDD.n233 20.5561
R4314 VDD.n231 VDD.n69 20.5561
R4315 VDD.n231 VDD.n230 20.5561
R4316 VDD.n236 VDD.n235 20.5561
R4317 VDD.n235 VDD.n234 20.5561
R4318 VDD.n220 VDD.n70 20.5561
R4319 VDD.n230 VDD.n70 20.5561
R4320 VDD.n269 VDD.n268 20.5561
R4321 VDD.n270 VDD.n269 20.5561
R4322 VDD.n256 VDD.n255 20.5561
R4323 VDD.n257 VDD.n256 20.5561
R4324 VDD.n272 VDD.n271 20.5561
R4325 VDD.n271 VDD.n270 20.5561
R4326 VDD.n240 VDD.n52 20.5561
R4327 VDD.n257 VDD.n52 20.5561
R4328 VDD.n19 VDD.n17 20.5561
R4329 VDD.n304 VDD.n19 20.5561
R4330 VDD.n290 VDD.n289 20.5561
R4331 VDD.n291 VDD.n290 20.5561
R4332 VDD.n26 VDD.n20 20.5561
R4333 VDD.n304 VDD.n20 20.5561
R4334 VDD.n293 VDD.n292 20.5561
R4335 VDD.n292 VDD.n291 20.5561
R4336 VDD.n372 VDD.n371 20.5561
R4337 VDD.n373 VDD.n372 20.5561
R4338 VDD.n364 VDD.n363 20.5561
R4339 VDD.n365 VDD.n364 20.5561
R4340 VDD.n375 VDD.n374 20.5561
R4341 VDD.n374 VDD.n373 20.5561
R4342 VDD.n317 VDD.n9 20.5561
R4343 VDD.n365 VDD.n9 20.5561
R4344 VDD.n350 VDD.n349 20.5561
R4345 VDD.n351 VDD.n350 20.5561
R4346 VDD.n353 VDD.n352 20.5561
R4347 VDD.n352 VDD.n351 20.5561
R4348 VDD.n354 VDD.n340 19.1
R4349 VDD.n125 VDD.n122 18.7082
R4350 VDD.n124 VDD.n123 18.7072
R4351 VDD.n492 VDD 18.0711
R4352 VDD.n495 VDD 18.0711
R4353 VDD.n531 VDD 18.0711
R4354 VDD.n534 VDD 18.0711
R4355 VDD.n570 VDD 18.0711
R4356 VDD.n573 VDD 18.0711
R4357 VDD.n609 VDD 18.0711
R4358 VDD.n612 VDD 18.0711
R4359 VDD.n990 VDD 18.0711
R4360 VDD.n987 VDD 18.0711
R4361 VDD.n961 VDD 18.0711
R4362 VDD.n958 VDD 18.0711
R4363 VDD.n932 VDD 18.0711
R4364 VDD.n929 VDD 18.0711
R4365 VDD.n903 VDD 18.0711
R4366 VDD.n900 VDD 18.0711
R4367 VDD.n874 VDD 18.0711
R4368 VDD.n871 VDD 18.0711
R4369 VDD.n845 VDD 18.0711
R4370 VDD.n842 VDD 18.0711
R4371 VDD.n816 VDD 18.0711
R4372 VDD.n443 VDD.t108 17.8272
R4373 VDD.n425 VDD.t165 17.8272
R4374 VDD.n407 VDD.t32 17.8272
R4375 VDD.n389 VDD.t42 17.8272
R4376 VDD.n994 VDD.t103 17.8272
R4377 VDD.n965 VDD.t114 17.8272
R4378 VDD.n936 VDD.t9 17.8272
R4379 VDD.n907 VDD.t166 17.8272
R4380 VDD.n878 VDD.t189 17.8272
R4381 VDD.n849 VDD.t85 17.8272
R4382 VDD.n820 VDD.t1 17.8272
R4383 VDD.n476 VDD.n475 17.7258
R4384 VDD.n515 VDD.n514 17.7258
R4385 VDD.n554 VDD.n553 17.7258
R4386 VDD.n593 VDD.n592 17.7258
R4387 VDD.n1004 VDD.n1003 17.7258
R4388 VDD.n975 VDD.n974 17.7258
R4389 VDD.n946 VDD.n945 17.7258
R4390 VDD.n917 VDD.n916 17.7258
R4391 VDD.n888 VDD.n887 17.7258
R4392 VDD.n859 VDD.n858 17.7258
R4393 VDD.n830 VDD.n829 17.7258
R4394 VDD.n118 VDD.n117 16.4845
R4395 VDD.n312 VDD.n311 16.4845
R4396 VDD.n39 VDD.n38 16.4845
R4397 VDD.n62 VDD.n61 16.4845
R4398 VDD.n184 VDD.n183 16.4845
R4399 VDD.n92 VDD.n91 16.4845
R4400 VDD.n331 VDD.t36 16.4465
R4401 VDD.n338 VDD.t138 16.4465
R4402 VDD.n162 VDD.t44 15.1423
R4403 VDD.n191 VDD.t136 15.1423
R4404 VDD.n86 VDD.t59 15.1423
R4405 VDD.n86 VDD.t52 15.1423
R4406 VDD.n188 VDD.t134 15.1423
R4407 VDD.n225 VDD.t112 15.1423
R4408 VDD.n225 VDD.t67 15.1423
R4409 VDD.n237 VDD.t30 15.1423
R4410 VDD.n51 VDD.t48 15.1423
R4411 VDD.n51 VDD.t183 15.1423
R4412 VDD.n277 VDD.t50 15.1423
R4413 VDD.n299 VDD.t69 15.1423
R4414 VDD.n299 VDD.t122 15.1423
R4415 VDD.n18 VDD.t91 15.1423
R4416 VDD.n8 VDD.t174 15.1423
R4417 VDD.n8 VDD.t18 15.1423
R4418 VDD.n376 VDD.t172 15.1423
R4419 VDD.n316 VDD.t164 15.1423
R4420 VDD.n295 VDD.t24 15.1423
R4421 VDD.n242 VDD.t61 15.1423
R4422 VDD.n222 VDD.t16 15.1423
R4423 VDD.n100 VDD.t5 15.1423
R4424 VDD.n165 VDD.t7 15.1423
R4425 VDD.n165 VDD.t3 15.1423
R4426 VDD.n32 VDD.n21 14.7003
R4427 VDD.n333 VDD.n329 14.6002
R4428 VDD.n334 VDD.n328 14.6002
R4429 VDD.n335 VDD.n327 14.6002
R4430 VDD.n336 VDD.n326 14.6002
R4431 VDD.n337 VDD.n325 14.6002
R4432 VDD.n141 VDD.n140 14.2846
R4433 VDD.n134 VDD.n132 13.357
R4434 VDD.n15 VDD.n11 13.2251
R4435 VDD.n287 VDD.n29 13.2251
R4436 VDD.n254 VDD.n54 13.2251
R4437 VDD.n181 VDD.n74 13.2251
R4438 VDD.n195 VDD.n90 13.2251
R4439 VDD.n154 VDD.n109 13.2251
R4440 VDD.n127 VDD.n126 13.0513
R4441 VDD.n477 VDD.n476 12.541
R4442 VDD.n516 VDD.n515 12.541
R4443 VDD.n555 VDD.n554 12.541
R4444 VDD.n594 VDD.n593 12.541
R4445 VDD.n1003 VDD.n1002 12.541
R4446 VDD.n974 VDD.n973 12.541
R4447 VDD.n945 VDD.n944 12.541
R4448 VDD.n916 VDD.n915 12.541
R4449 VDD.n887 VDD.n886 12.541
R4450 VDD.n858 VDD.n857 12.541
R4451 VDD.n829 VDD.n828 12.541
R4452 VDD.n273 VDD.n44 12.4146
R4453 VDD.n154 VDD.t63 11.9046
R4454 VDD.n178 VDD.t170 11.9046
R4455 VDD.n195 VDD.t178 11.9046
R4456 VDD.n82 VDD.t118 11.9046
R4457 VDD.n247 VDD.t144 11.9046
R4458 VDD.n281 VDD.t71 11.9046
R4459 VDD.n309 VDD.t227 11.9046
R4460 VDD.n148 VDD.t83 11.9046
R4461 VDD.n11 VDD.t231 11.9046
R4462 VDD.n287 VDD.t22 11.9046
R4463 VDD.n254 VDD.t146 11.9046
R4464 VDD.n181 VDD.t120 11.9046
R4465 VDD.n285 VDD.n21 11.2431
R4466 VDD.n309 VDD.n308 11.2069
R4467 VDD.n247 VDD.n60 11.2069
R4468 VDD.n187 VDD.n82 11.2069
R4469 VDD.n178 VDD.n95 11.2069
R4470 VDD.n126 VDD.n120 11.1021
R4471 VDD.n116 VDD.n113 10.8829
R4472 VDD.n150 VDD.n113 10.8829
R4473 VDD.n114 VDD.n110 10.8829
R4474 VDD.n150 VDD.n114 10.8829
R4475 VDD.n96 VDD.n80 10.8829
R4476 VDD.n175 VDD.n96 10.8829
R4477 VDD.n101 VDD.n97 10.8829
R4478 VDD.n175 VDD.n97 10.8829
R4479 VDD.n216 VDD.n215 10.8829
R4480 VDD.n217 VDD.n216 10.8829
R4481 VDD.n219 VDD.n218 10.8829
R4482 VDD.n218 VDD.n217 10.8829
R4483 VDD.n56 VDD.n49 10.8829
R4484 VDD.n250 VDD.n56 10.8829
R4485 VDD.n239 VDD.n57 10.8829
R4486 VDD.n250 VDD.n57 10.8829
R4487 VDD.n265 VDD.n34 10.8829
R4488 VDD.n284 VDD.n34 10.8829
R4489 VDD.n35 VDD.n30 10.8829
R4490 VDD.n284 VDD.n35 10.8829
R4491 VDD.n361 VDD.n360 10.8829
R4492 VDD.n360 VDD.n359 10.8829
R4493 VDD.n320 VDD.n319 10.8829
R4494 VDD.n359 VDD.n320 10.8829
R4495 VDD.n266 VDD 10.4678
R4496 VDD.n44 VDD.n43 10.1531
R4497 VDD.n281 VDD.n37 10.0007
R4498 VDD.n479 VDD.n449 9.5406
R4499 VDD.n518 VDD.n431 9.5406
R4500 VDD.n557 VDD.n413 9.5406
R4501 VDD.n596 VDD.n395 9.5406
R4502 VDD.n633 VDD.n631 9.5406
R4503 VDD.n661 VDD.n659 9.5406
R4504 VDD.n689 VDD.n687 9.5406
R4505 VDD.n717 VDD.n715 9.5406
R4506 VDD.n745 VDD.n743 9.5406
R4507 VDD.n773 VDD.n771 9.5406
R4508 VDD.n801 VDD.n799 9.5406
R4509 VDD VDD.n457 9.3245
R4510 VDD.n614 VDD.n387 9.3005
R4511 VDD.n605 VDD.n604 9.3005
R4512 VDD.n606 VDD.n605 9.3005
R4513 VDD.n596 VDD.n595 9.3005
R4514 VDD.n597 VDD.n596 9.3005
R4515 VDD.n575 VDD.n405 9.3005
R4516 VDD.n578 VDD.n577 9.3005
R4517 VDD.n581 VDD.n580 9.3005
R4518 VDD.n566 VDD.n565 9.3005
R4519 VDD.n567 VDD.n566 9.3005
R4520 VDD.n557 VDD.n556 9.3005
R4521 VDD.n558 VDD.n557 9.3005
R4522 VDD.n536 VDD.n423 9.3005
R4523 VDD.n539 VDD.n538 9.3005
R4524 VDD.n542 VDD.n541 9.3005
R4525 VDD.n527 VDD.n526 9.3005
R4526 VDD.n528 VDD.n527 9.3005
R4527 VDD.n518 VDD.n517 9.3005
R4528 VDD.n519 VDD.n518 9.3005
R4529 VDD.n497 VDD.n441 9.3005
R4530 VDD.n500 VDD.n499 9.3005
R4531 VDD.n503 VDD.n502 9.3005
R4532 VDD.n488 VDD.n487 9.3005
R4533 VDD.n489 VDD.n488 9.3005
R4534 VDD.n479 VDD.n478 9.3005
R4535 VDD.n480 VDD.n479 9.3005
R4536 VDD.n458 VDD.n456 9.3005
R4537 VDD.n461 VDD.n460 9.3005
R4538 VDD.n464 VDD.n463 9.3005
R4539 VDD.n615 VDD.n385 9.3005
R4540 VDD.n613 VDD.n612 9.3005
R4541 VDD.n609 VDD.n608 9.3005
R4542 VDD.n607 VDD.n388 9.3005
R4543 VDD.n603 VDD.n602 9.3005
R4544 VDD.n599 VDD.n598 9.3005
R4545 VDD.n394 VDD.n391 9.3005
R4546 VDD.n591 VDD.n590 9.3005
R4547 VDD.n589 VDD.n588 9.3005
R4548 VDD.n404 VDD.n396 9.3005
R4549 VDD.n583 VDD.n582 9.3005
R4550 VDD.n576 VDD.n403 9.3005
R4551 VDD.n574 VDD.n573 9.3005
R4552 VDD.n570 VDD.n569 9.3005
R4553 VDD.n568 VDD.n406 9.3005
R4554 VDD.n564 VDD.n563 9.3005
R4555 VDD.n560 VDD.n559 9.3005
R4556 VDD.n412 VDD.n409 9.3005
R4557 VDD.n552 VDD.n551 9.3005
R4558 VDD.n550 VDD.n549 9.3005
R4559 VDD.n422 VDD.n414 9.3005
R4560 VDD.n544 VDD.n543 9.3005
R4561 VDD.n537 VDD.n421 9.3005
R4562 VDD.n535 VDD.n534 9.3005
R4563 VDD.n531 VDD.n530 9.3005
R4564 VDD.n529 VDD.n424 9.3005
R4565 VDD.n525 VDD.n524 9.3005
R4566 VDD.n521 VDD.n520 9.3005
R4567 VDD.n430 VDD.n427 9.3005
R4568 VDD.n513 VDD.n512 9.3005
R4569 VDD.n511 VDD.n510 9.3005
R4570 VDD.n440 VDD.n432 9.3005
R4571 VDD.n505 VDD.n504 9.3005
R4572 VDD.n498 VDD.n439 9.3005
R4573 VDD.n496 VDD.n495 9.3005
R4574 VDD.n492 VDD.n491 9.3005
R4575 VDD.n490 VDD.n442 9.3005
R4576 VDD.n486 VDD.n485 9.3005
R4577 VDD.n482 VDD.n481 9.3005
R4578 VDD.n448 VDD.n445 9.3005
R4579 VDD.n474 VDD.n473 9.3005
R4580 VDD.n472 VDD.n471 9.3005
R4581 VDD.n455 VDD.n450 9.3005
R4582 VDD.n466 VDD.n465 9.3005
R4583 VDD.n459 VDD.n454 9.3005
R4584 VDD.n823 VDD.n822 9.3005
R4585 VDD.n822 VDD.n819 9.3005
R4586 VDD.n801 VDD.n800 9.3005
R4587 VDD.n802 VDD.n801 9.3005
R4588 VDD.n786 VDD.n785 9.3005
R4589 VDD.n839 VDD.n838 9.3005
R4590 VDD.n836 VDD.n835 9.3005
R4591 VDD.n852 VDD.n851 9.3005
R4592 VDD.n851 VDD.n848 9.3005
R4593 VDD.n773 VDD.n772 9.3005
R4594 VDD.n774 VDD.n773 9.3005
R4595 VDD.n758 VDD.n757 9.3005
R4596 VDD.n868 VDD.n867 9.3005
R4597 VDD.n865 VDD.n864 9.3005
R4598 VDD.n881 VDD.n880 9.3005
R4599 VDD.n880 VDD.n877 9.3005
R4600 VDD.n745 VDD.n744 9.3005
R4601 VDD.n746 VDD.n745 9.3005
R4602 VDD.n730 VDD.n729 9.3005
R4603 VDD.n897 VDD.n896 9.3005
R4604 VDD.n894 VDD.n893 9.3005
R4605 VDD.n910 VDD.n909 9.3005
R4606 VDD.n909 VDD.n906 9.3005
R4607 VDD.n717 VDD.n716 9.3005
R4608 VDD.n718 VDD.n717 9.3005
R4609 VDD.n702 VDD.n701 9.3005
R4610 VDD.n926 VDD.n925 9.3005
R4611 VDD.n923 VDD.n922 9.3005
R4612 VDD.n939 VDD.n938 9.3005
R4613 VDD.n938 VDD.n935 9.3005
R4614 VDD.n689 VDD.n688 9.3005
R4615 VDD.n690 VDD.n689 9.3005
R4616 VDD.n674 VDD.n673 9.3005
R4617 VDD.n955 VDD.n954 9.3005
R4618 VDD.n952 VDD.n951 9.3005
R4619 VDD.n968 VDD.n967 9.3005
R4620 VDD.n967 VDD.n964 9.3005
R4621 VDD.n661 VDD.n660 9.3005
R4622 VDD.n662 VDD.n661 9.3005
R4623 VDD.n646 VDD.n645 9.3005
R4624 VDD.n984 VDD.n983 9.3005
R4625 VDD.n981 VDD.n980 9.3005
R4626 VDD.n997 VDD.n996 9.3005
R4627 VDD.n996 VDD.n993 9.3005
R4628 VDD.n633 VDD.n632 9.3005
R4629 VDD.n634 VDD.n633 9.3005
R4630 VDD.n816 VDD.n815 9.3005
R4631 VDD.n818 VDD.n817 9.3005
R4632 VDD.n807 VDD.n806 9.3005
R4633 VDD.n825 VDD.n824 9.3005
R4634 VDD.n827 VDD.n826 9.3005
R4635 VDD.n803 VDD.n798 9.3005
R4636 VDD.n832 VDD.n831 9.3005
R4637 VDD.n834 VDD.n833 9.3005
R4638 VDD.n787 VDD.n784 9.3005
R4639 VDD.n841 VDD.n840 9.3005
R4640 VDD.n843 VDD.n842 9.3005
R4641 VDD.n845 VDD.n844 9.3005
R4642 VDD.n847 VDD.n846 9.3005
R4643 VDD.n779 VDD.n778 9.3005
R4644 VDD.n854 VDD.n853 9.3005
R4645 VDD.n856 VDD.n855 9.3005
R4646 VDD.n775 VDD.n770 9.3005
R4647 VDD.n861 VDD.n860 9.3005
R4648 VDD.n863 VDD.n862 9.3005
R4649 VDD.n759 VDD.n756 9.3005
R4650 VDD.n870 VDD.n869 9.3005
R4651 VDD.n872 VDD.n871 9.3005
R4652 VDD.n874 VDD.n873 9.3005
R4653 VDD.n876 VDD.n875 9.3005
R4654 VDD.n751 VDD.n750 9.3005
R4655 VDD.n883 VDD.n882 9.3005
R4656 VDD.n885 VDD.n884 9.3005
R4657 VDD.n747 VDD.n742 9.3005
R4658 VDD.n890 VDD.n889 9.3005
R4659 VDD.n892 VDD.n891 9.3005
R4660 VDD.n731 VDD.n728 9.3005
R4661 VDD.n899 VDD.n898 9.3005
R4662 VDD.n901 VDD.n900 9.3005
R4663 VDD.n903 VDD.n902 9.3005
R4664 VDD.n905 VDD.n904 9.3005
R4665 VDD.n723 VDD.n722 9.3005
R4666 VDD.n912 VDD.n911 9.3005
R4667 VDD.n914 VDD.n913 9.3005
R4668 VDD.n719 VDD.n714 9.3005
R4669 VDD.n919 VDD.n918 9.3005
R4670 VDD.n921 VDD.n920 9.3005
R4671 VDD.n703 VDD.n700 9.3005
R4672 VDD.n928 VDD.n927 9.3005
R4673 VDD.n930 VDD.n929 9.3005
R4674 VDD.n932 VDD.n931 9.3005
R4675 VDD.n934 VDD.n933 9.3005
R4676 VDD.n695 VDD.n694 9.3005
R4677 VDD.n941 VDD.n940 9.3005
R4678 VDD.n943 VDD.n942 9.3005
R4679 VDD.n691 VDD.n686 9.3005
R4680 VDD.n948 VDD.n947 9.3005
R4681 VDD.n950 VDD.n949 9.3005
R4682 VDD.n675 VDD.n672 9.3005
R4683 VDD.n957 VDD.n956 9.3005
R4684 VDD.n959 VDD.n958 9.3005
R4685 VDD.n961 VDD.n960 9.3005
R4686 VDD.n963 VDD.n962 9.3005
R4687 VDD.n667 VDD.n666 9.3005
R4688 VDD.n970 VDD.n969 9.3005
R4689 VDD.n972 VDD.n971 9.3005
R4690 VDD.n663 VDD.n658 9.3005
R4691 VDD.n977 VDD.n976 9.3005
R4692 VDD.n979 VDD.n978 9.3005
R4693 VDD.n647 VDD.n644 9.3005
R4694 VDD.n986 VDD.n985 9.3005
R4695 VDD.n988 VDD.n987 9.3005
R4696 VDD.n990 VDD.n989 9.3005
R4697 VDD.n992 VDD.n991 9.3005
R4698 VDD.n639 VDD.n638 9.3005
R4699 VDD.n999 VDD.n998 9.3005
R4700 VDD.n1001 VDD.n1000 9.3005
R4701 VDD.n635 VDD.n630 9.3005
R4702 VDD.n618 VDD.n617 9.3005
R4703 VDD.n621 VDD.n620 9.3005
R4704 VDD.n629 VDD.n628 9.3005
R4705 VDD.n386 VDD.n378 9.3005
R4706 VDD.n623 VDD.n622 9.3005
R4707 VDD.n268 VDD.n267 8.39406
R4708 VDD.n42 VDD.n41 7.40898
R4709 VDD.n449 VDD 7.01471
R4710 VDD.n431 VDD 7.01471
R4711 VDD.n413 VDD 7.01471
R4712 VDD.n395 VDD 7.01471
R4713 VDD.n631 VDD 7.01471
R4714 VDD.n659 VDD 7.01471
R4715 VDD.n687 VDD 7.01471
R4716 VDD.n715 VDD 7.01471
R4717 VDD.n743 VDD 7.01471
R4718 VDD.n771 VDD 7.01471
R4719 VDD.n799 VDD 7.01471
R4720 VDD.n371 VDD.n370 6.79942
R4721 VDD.n289 VDD.n288 6.74738
R4722 VDD.n255 VDD.n50 6.74738
R4723 VDD.n228 VDD.n69 6.74738
R4724 VDD.n201 VDD.n200 6.74738
R4725 VDD.n156 VDD.n155 6.74738
R4726 VDD.n276 VDD.n43 6.54595
R4727 VDD.n303 VDD.n302 6.48514
R4728 VDD.n42 VDD.n37 6.43879
R4729 VDD.n268 VDD.n263 6.43519
R4730 VDD.n264 VDD.n17 6.14034
R4731 VDD.n72 VDD.n59 6.14034
R4732 VDD.n214 VDD.n213 6.14034
R4733 VDD.n115 VDD.n94 6.14034
R4734 VDD.n118 VDD.n112 5.88536
R4735 VDD.n313 VDD.n312 5.88536
R4736 VDD.n39 VDD.n33 5.88536
R4737 VDD.n62 VDD.n55 5.88536
R4738 VDD.n184 VDD.n182 5.88536
R4739 VDD.n194 VDD.n92 5.88536
R4740 VDD.n147 VDD.n118 5.86002
R4741 VDD.n312 VDD.n310 5.86002
R4742 VDD.n280 VDD.n39 5.86002
R4743 VDD.n246 VDD.n62 5.86002
R4744 VDD.n185 VDD.n184 5.86002
R4745 VDD.n179 VDD.n92 5.86002
R4746 VDD.n363 VDD.n362 5.75877
R4747 VDD.n133 VDD.n128 4.42757
R4748 VDD.n461 VDD.n456 4.36685
R4749 VDD.n500 VDD.n441 4.36685
R4750 VDD.n539 VDD.n423 4.36685
R4751 VDD.n578 VDD.n405 4.36685
R4752 VDD.n618 VDD.n387 4.36685
R4753 VDD.n983 VDD.n646 4.36685
R4754 VDD.n954 VDD.n674 4.36685
R4755 VDD.n925 VDD.n702 4.36685
R4756 VDD.n896 VDD.n730 4.36685
R4757 VDD.n867 VDD.n758 4.36685
R4758 VDD.n838 VDD.n786 4.36685
R4759 VDD.n111 VDD.n109 3.93667
R4760 VDD.n151 VDD.n111 3.93667
R4761 VDD.n167 VDD.n166 3.93667
R4762 VDD.n168 VDD.n167 3.93667
R4763 VDD.n171 VDD.n95 3.93667
R4764 VDD.n172 VDD.n171 3.93667
R4765 VDD.n90 VDD.n88 3.93667
R4766 VDD.n173 VDD.n88 3.93667
R4767 VDD.n197 VDD.n196 3.93667
R4768 VDD.n198 VDD.n197 3.93667
R4769 VDD.n187 VDD.n84 3.93667
R4770 VDD.n210 VDD.n84 3.93667
R4771 VDD.n74 VDD.n68 3.93667
R4772 VDD.n78 VDD.n68 3.93667
R4773 VDD.n226 VDD.n67 3.93667
R4774 VDD.n71 VDD.n67 3.93667
R4775 VDD.n66 VDD.n60 3.93667
R4776 VDD.n66 VDD.n58 3.93667
R4777 VDD.n54 VDD.n53 3.93667
R4778 VDD.n251 VDD.n53 3.93667
R4779 VDD.n261 VDD.n260 3.93667
R4780 VDD.n260 VDD.n259 3.93667
R4781 VDD.n47 VDD.n41 3.93667
R4782 VDD.n47 VDD.n36 3.93667
R4783 VDD.n31 VDD.n29 3.93667
R4784 VDD.n32 VDD.n31 3.93667
R4785 VDD.n301 VDD.n300 3.93667
R4786 VDD.n302 VDD.n301 3.93667
R4787 VDD.n308 VDD.n307 3.93667
R4788 VDD.n307 VDD.n306 3.93667
R4789 VDD.n15 VDD.n10 3.93667
R4790 VDD.n321 VDD.n10 3.93667
R4791 VDD.n369 VDD.n368 3.93667
R4792 VDD.n368 VDD.n367 3.93667
R4793 VDD.n5 VDD.n2 3.93667
R4794 VDD.n356 VDD.n355 3.93667
R4795 VDD.n357 VDD.n356 3.93667
R4796 VDD.n342 VDD.n322 3.93667
R4797 VDD.n357 VDD.n322 3.93667
R4798 VDD.n341 VDD.n323 3.85467
R4799 VDD.n343 VDD.n324 3.85467
R4800 VDD.n142 VDD.n121 3.75923
R4801 VDD.n444 VDD 3.7406
R4802 VDD.n426 VDD 3.7406
R4803 VDD.n408 VDD 3.7406
R4804 VDD.n390 VDD 3.7406
R4805 VDD.n995 VDD 3.7406
R4806 VDD.n966 VDD 3.7406
R4807 VDD.n937 VDD 3.7406
R4808 VDD.n908 VDD 3.7406
R4809 VDD.n879 VDD 3.7406
R4810 VDD.n850 VDD 3.7406
R4811 VDD.n821 VDD 3.7406
R4812 VDD.n149 VDD.n148 3.08383
R4813 VDD.n154 VDD.n153 3.08383
R4814 VDD.n153 VDD.n152 3.08383
R4815 VDD.n178 VDD.n177 3.08383
R4816 VDD.n177 VDD.n176 3.08383
R4817 VDD.n195 VDD.n89 3.08383
R4818 VDD.n174 VDD.n89 3.08383
R4819 VDD.n82 VDD.n76 3.08383
R4820 VDD.n209 VDD.n76 3.08383
R4821 VDD.n181 VDD.n77 3.08383
R4822 VDD.n79 VDD.n77 3.08383
R4823 VDD.n248 VDD.n247 3.08383
R4824 VDD.n249 VDD.n248 3.08383
R4825 VDD.n254 VDD.n253 3.08383
R4826 VDD.n253 VDD.n252 3.08383
R4827 VDD.n282 VDD.n281 3.08383
R4828 VDD.n283 VDD.n282 3.08383
R4829 VDD.n287 VDD.n286 3.08383
R4830 VDD.n286 VDD.n285 3.08383
R4831 VDD.n309 VDD.n12 3.08383
R4832 VDD.n305 VDD.n12 3.08383
R4833 VDD.n13 VDD.n11 3.08383
R4834 VDD.n358 VDD.n13 3.08383
R4835 VDD.n274 VDD.n273 2.84494
R4836 VDD.n462 VDD.n461 2.81171
R4837 VDD.n501 VDD.n500 2.81171
R4838 VDD.n540 VDD.n539 2.81171
R4839 VDD.n579 VDD.n578 2.81171
R4840 VDD.n619 VDD.n618 2.81171
R4841 VDD.n983 VDD.n982 2.81171
R4842 VDD.n954 VDD.n953 2.81171
R4843 VDD.n925 VDD.n924 2.81171
R4844 VDD.n896 VDD.n895 2.81171
R4845 VDD.n867 VDD.n866 2.81171
R4846 VDD.n838 VDD.n837 2.81171
R4847 VDD.n376 VDD.n2 2.74336
R4848 VDD.n358 VDD.n357 2.59436
R4849 VDD.n463 VDD.n462 2.45284
R4850 VDD.n502 VDD.n501 2.45284
R4851 VDD.n541 VDD.n540 2.45284
R4852 VDD.n580 VDD.n579 2.45284
R4853 VDD.n620 VDD.n619 2.45284
R4854 VDD.n982 VDD.n981 2.45284
R4855 VDD.n953 VDD.n952 2.45284
R4856 VDD.n924 VDD.n923 2.45284
R4857 VDD.n895 VDD.n894 2.45284
R4858 VDD.n866 VDD.n865 2.45284
R4859 VDD.n837 VDD.n836 2.45284
R4860 VDD.n329 VDD.t140 1.84683
R4861 VDD.n329 VDD.t142 1.84683
R4862 VDD.n328 VDD.t75 1.84683
R4863 VDD.n328 VDD.t132 1.84683
R4864 VDD.n327 VDD.t38 1.84683
R4865 VDD.n327 VDD.t40 1.84683
R4866 VDD.n326 VDD.t77 1.84683
R4867 VDD.n326 VDD.t79 1.84683
R4868 VDD.n325 VDD.t185 1.84683
R4869 VDD.n325 VDD.t187 1.84683
R4870 VDD.n369 VDD.n8 1.52129
R4871 VDD.n300 VDD.n299 1.52129
R4872 VDD.n261 VDD.n51 1.52129
R4873 VDD.n226 VDD.n225 1.52129
R4874 VDD.n196 VDD.n86 1.52129
R4875 VDD.n166 VDD.n165 1.52129
R4876 VDD.n155 VDD.n104 1.46295
R4877 VDD.n200 VDD.n199 1.46295
R4878 VDD.n229 VDD.n228 1.46295
R4879 VDD.n258 VDD.n50 1.46295
R4880 VDD.n288 VDD.n22 1.46295
R4881 VDD.n366 VDD.n7 1.46295
R4882 VDD.n117 VDD.t34 1.45813
R4883 VDD.n117 VDD.t65 1.45813
R4884 VDD.n311 VDD.t233 1.45813
R4885 VDD.n311 VDD.t229 1.45813
R4886 VDD.n38 VDD.t73 1.45813
R4887 VDD.n38 VDD.t20 1.45813
R4888 VDD.n61 VDD.t26 1.45813
R4889 VDD.n61 VDD.t28 1.45813
R4890 VDD.n183 VDD.t150 1.45813
R4891 VDD.n183 VDD.t148 1.45813
R4892 VDD.n91 VDD.t168 1.45813
R4893 VDD.n91 VDD.t176 1.45813
R4894 VDD.n277 VDD.n41 1.39686
R4895 VDD.n316 VDD.n15 1.09244
R4896 VDD.n295 VDD.n29 1.09244
R4897 VDD.n242 VDD.n54 1.09244
R4898 VDD.n222 VDD.n74 1.09244
R4899 VDD.n191 VDD.n90 1.09244
R4900 VDD.n162 VDD.n109 1.09244
R4901 VDD.n362 VDD.n7 0.989118
R4902 VDD.n147 VDD.n146 0.988365
R4903 VDD.n310 VDD.n16 0.988365
R4904 VDD.n280 VDD.n279 0.988365
R4905 VDD.n246 VDD.n245 0.988365
R4906 VDD.n186 VDD.n185 0.988365
R4907 VDD.n180 VDD.n179 0.988365
R4908 VDD.n112 VDD.n108 0.984009
R4909 VDD.n314 VDD.n313 0.984009
R4910 VDD.n33 VDD.n28 0.984009
R4911 VDD.n244 VDD.n55 0.984009
R4912 VDD.n182 VDD.n73 0.984009
R4913 VDD.n194 VDD.n193 0.984009
R4914 VDD.n144 VDD.n143 0.972503
R4915 VDD.n308 VDD.n18 0.925801
R4916 VDD.n237 VDD.n60 0.925801
R4917 VDD.n188 VDD.n187 0.925801
R4918 VDD.n100 VDD.n95 0.925801
R4919 VDD.n163 VDD.n162 0.921929
R4920 VDD.n192 VDD.n191 0.921929
R4921 VDD.n316 VDD.n315 0.921929
R4922 VDD.n296 VDD.n295 0.921929
R4923 VDD.n243 VDD.n242 0.921929
R4924 VDD.n223 VDD.n222 0.921929
R4925 VDD.n189 VDD.n188 0.908023
R4926 VDD.n237 VDD.n63 0.908023
R4927 VDD.n278 VDD.n277 0.908023
R4928 VDD.n297 VDD.n18 0.908023
R4929 VDD.n377 VDD.n376 0.908023
R4930 VDD.n100 VDD.n93 0.908023
R4931 VDD.n475 VDD 0.755
R4932 VDD.n514 VDD 0.755
R4933 VDD.n553 VDD 0.755
R4934 VDD.n592 VDD 0.755
R4935 VDD VDD.n975 0.755
R4936 VDD VDD.n946 0.755
R4937 VDD VDD.n917 0.755
R4938 VDD VDD.n888 0.755
R4939 VDD VDD.n859 0.755
R4940 VDD VDD.n830 0.755
R4941 VDD.n275 VDD.n44 0.682885
R4942 VDD.n264 VDD.n25 0.659579
R4943 VDD.n227 VDD.n72 0.659579
R4944 VDD.n214 VDD.n81 0.659579
R4945 VDD.n115 VDD.n106 0.659579
R4946 VDD.n168 VDD.n104 0.649112
R4947 VDD.n199 VDD.n198 0.649112
R4948 VDD.n229 VDD.n71 0.649112
R4949 VDD.n259 VDD.n258 0.649112
R4950 VDD.n302 VDD.n22 0.648964
R4951 VDD.n367 VDD.n366 0.648964
R4952 VDD.n339 VDD.n338 0.643506
R4953 VDD.n1005 VDD 0.6255
R4954 VDD.n344 VDD.n0 0.610727
R4955 VDD.n140 VDD.n139 0.601149
R4956 VDD.n139 VDD.n138 0.601149
R4957 VDD.n135 VDD.n134 0.601149
R4958 VDD.n136 VDD.n135 0.601149
R4959 VDD VDD.n1007 0.553005
R4960 VDD.n133 VDD.n130 0.405314
R4961 VDD.n137 VDD.n130 0.405314
R4962 VDD.n129 VDD.n121 0.405314
R4963 VDD.n131 VDD.n129 0.405314
R4964 VDD.n814 VDD 0.385917
R4965 VDD.n814 VDD 0.385917
R4966 VDD.n263 VDD.n262 0.364728
R4967 VDD.n1005 VDD.n1004 0.359
R4968 VDD.n126 VDD 0.331269
R4969 VDD.n190 VDD.n86 0.317443
R4970 VDD.n225 VDD.n224 0.317443
R4971 VDD.n51 VDD.n40 0.317443
R4972 VDD.n299 VDD.n298 0.317443
R4973 VDD.n8 VDD.n1 0.317443
R4974 VDD.n165 VDD.n164 0.317443
R4975 VDD.n1007 VDD.n1006 0.279456
R4976 VDD.n1006 VDD.n1005 0.27291
R4977 VDD.n814 VDD 0.240083
R4978 VDD.n148 VDD.n147 0.179346
R4979 VDD.n313 VDD.n11 0.179346
R4980 VDD.n310 VDD.n309 0.179346
R4981 VDD.n287 VDD.n33 0.179346
R4982 VDD.n281 VDD.n280 0.179346
R4983 VDD.n254 VDD.n55 0.179346
R4984 VDD.n247 VDD.n246 0.179346
R4985 VDD.n182 VDD.n181 0.179346
R4986 VDD.n185 VDD.n82 0.179346
R4987 VDD.n195 VDD.n194 0.179346
R4988 VDD.n179 VDD.n178 0.179346
R4989 VDD.n154 VDD.n112 0.179346
R4990 VDD.n145 VDD.n144 0.158248
R4991 VDD.n1006 VDD 0.122512
R4992 VDD.n338 VDD.n337 0.0814285
R4993 VDD.n337 VDD.n336 0.0814285
R4994 VDD.n336 VDD.n335 0.0814285
R4995 VDD.n335 VDD.n334 0.0814285
R4996 VDD.n334 VDD.n333 0.0814285
R4997 VDD.n124 VDD 0.0649231
R4998 VDD VDD.n125 0.0639615
R4999 VDD.n123 VDD 0.063
R5000 VDD.n122 VDD 0.063
R5001 VDD.n488 VDD.n444 0.057952
R5002 VDD.n527 VDD.n426 0.057952
R5003 VDD.n566 VDD.n408 0.057952
R5004 VDD.n605 VDD.n390 0.057952
R5005 VDD.n996 VDD.n995 0.057952
R5006 VDD.n967 VDD.n966 0.057952
R5007 VDD.n938 VDD.n937 0.057952
R5008 VDD.n909 VDD.n908 0.057952
R5009 VDD.n880 VDD.n879 0.057952
R5010 VDD.n851 VDD.n850 0.057952
R5011 VDD.n822 VDD.n821 0.057952
R5012 VDD.n370 VDD.n7 0.0525325
R5013 VDD.n288 VDD.n25 0.0525325
R5014 VDD.n262 VDD.n50 0.0525325
R5015 VDD.n228 VDD.n227 0.0525325
R5016 VDD.n200 VDD.n81 0.0525325
R5017 VDD.n155 VDD.n106 0.0525325
R5018 VDD.n146 VDD.n145 0.0492521
R5019 VDD.n146 VDD.n108 0.0485075
R5020 VDD.n193 VDD.n180 0.0485075
R5021 VDD.n186 VDD.n73 0.0485075
R5022 VDD.n245 VDD.n244 0.0485075
R5023 VDD.n279 VDD.n28 0.0485075
R5024 VDD.n314 VDD.n16 0.0485075
R5025 VDD.n332 VDD.n331 0.0419053
R5026 VDD.n333 VDD.n332 0.0400232
R5027 VDD.n491 VDD 0.04
R5028 VDD.n530 VDD 0.04
R5029 VDD.n569 VDD 0.04
R5030 VDD.n608 VDD 0.04
R5031 VDD.n989 VDD 0.04
R5032 VDD.n960 VDD 0.04
R5033 VDD.n931 VDD 0.04
R5034 VDD.n902 VDD 0.04
R5035 VDD.n873 VDD 0.04
R5036 VDD.n844 VDD 0.04
R5037 VDD.n815 VDD 0.04
R5038 VDD.n1007 VDD.n377 0.037294
R5039 VDD.n487 VDD 0.0365
R5040 VDD.n526 VDD 0.0365
R5041 VDD.n565 VDD 0.0365
R5042 VDD.n604 VDD 0.0365
R5043 VDD VDD.n997 0.0365
R5044 VDD VDD.n968 0.0365
R5045 VDD VDD.n939 0.0365
R5046 VDD VDD.n910 0.0365
R5047 VDD VDD.n881 0.0365
R5048 VDD VDD.n852 0.0365
R5049 VDD VDD.n823 0.0365
R5050 VDD.n132 VDD.n119 0.0332465
R5051 VDD.n141 VDD.n120 0.0332465
R5052 VDD.n331 VDD.n0 0.0323381
R5053 VDD.n481 VDD 0.032
R5054 VDD.n520 VDD 0.032
R5055 VDD.n559 VDD 0.032
R5056 VDD.n598 VDD 0.032
R5057 VDD.n998 VDD 0.032
R5058 VDD.n969 VDD 0.032
R5059 VDD.n940 VDD 0.032
R5060 VDD.n911 VDD 0.032
R5061 VDD.n882 VDD 0.032
R5062 VDD.n853 VDD 0.032
R5063 VDD.n824 VDD 0.032
R5064 VDD.n164 VDD.n93 0.0305923
R5065 VDD.n190 VDD.n189 0.0305923
R5066 VDD.n224 VDD.n63 0.0305923
R5067 VDD.n278 VDD.n40 0.0305923
R5068 VDD.n298 VDD.n297 0.0305923
R5069 VDD.n377 VDD.n1 0.0305923
R5070 VDD.n164 VDD.n163 0.0298914
R5071 VDD.n192 VDD.n190 0.0298914
R5072 VDD.n224 VDD.n223 0.0298914
R5073 VDD.n243 VDD.n40 0.0298914
R5074 VDD.n298 VDD.n296 0.0298914
R5075 VDD.n315 VDD.n1 0.0298914
R5076 VDD.n465 VDD 0.0245
R5077 VDD VDD.n455 0.0245
R5078 VDD.n455 VDD 0.0245
R5079 VDD.n472 VDD 0.0245
R5080 VDD.n489 VDD 0.0245
R5081 VDD.n496 VDD 0.0245
R5082 VDD VDD.n496 0.0245
R5083 VDD.n504 VDD 0.0245
R5084 VDD VDD.n440 0.0245
R5085 VDD.n440 VDD 0.0245
R5086 VDD.n511 VDD 0.0245
R5087 VDD.n528 VDD 0.0245
R5088 VDD.n535 VDD 0.0245
R5089 VDD VDD.n535 0.0245
R5090 VDD.n543 VDD 0.0245
R5091 VDD VDD.n422 0.0245
R5092 VDD.n422 VDD 0.0245
R5093 VDD.n550 VDD 0.0245
R5094 VDD.n567 VDD 0.0245
R5095 VDD.n574 VDD 0.0245
R5096 VDD VDD.n574 0.0245
R5097 VDD.n582 VDD 0.0245
R5098 VDD VDD.n404 0.0245
R5099 VDD.n404 VDD 0.0245
R5100 VDD.n589 VDD 0.0245
R5101 VDD.n606 VDD 0.0245
R5102 VDD.n613 VDD 0.0245
R5103 VDD VDD.n613 0.0245
R5104 VDD.n993 VDD 0.0245
R5105 VDD VDD.n988 0.0245
R5106 VDD.n988 VDD 0.0245
R5107 VDD.n647 VDD 0.0245
R5108 VDD VDD.n979 0.0245
R5109 VDD.n979 VDD 0.0245
R5110 VDD.n976 VDD 0.0245
R5111 VDD.n964 VDD 0.0245
R5112 VDD VDD.n959 0.0245
R5113 VDD.n959 VDD 0.0245
R5114 VDD.n675 VDD 0.0245
R5115 VDD VDD.n950 0.0245
R5116 VDD.n950 VDD 0.0245
R5117 VDD.n947 VDD 0.0245
R5118 VDD.n935 VDD 0.0245
R5119 VDD VDD.n930 0.0245
R5120 VDD.n930 VDD 0.0245
R5121 VDD.n703 VDD 0.0245
R5122 VDD VDD.n921 0.0245
R5123 VDD.n921 VDD 0.0245
R5124 VDD.n918 VDD 0.0245
R5125 VDD.n906 VDD 0.0245
R5126 VDD VDD.n901 0.0245
R5127 VDD.n901 VDD 0.0245
R5128 VDD.n731 VDD 0.0245
R5129 VDD VDD.n892 0.0245
R5130 VDD.n892 VDD 0.0245
R5131 VDD.n889 VDD 0.0245
R5132 VDD.n877 VDD 0.0245
R5133 VDD VDD.n872 0.0245
R5134 VDD.n872 VDD 0.0245
R5135 VDD.n759 VDD 0.0245
R5136 VDD VDD.n863 0.0245
R5137 VDD.n863 VDD 0.0245
R5138 VDD.n860 VDD 0.0245
R5139 VDD.n848 VDD 0.0245
R5140 VDD VDD.n843 0.0245
R5141 VDD.n843 VDD 0.0245
R5142 VDD.n787 VDD 0.0245
R5143 VDD VDD.n834 0.0245
R5144 VDD.n834 VDD 0.0245
R5145 VDD.n831 VDD 0.0245
R5146 VDD.n819 VDD 0.0245
R5147 VDD.n622 VDD 0.0244044
R5148 VDD VDD.n386 0.0244044
R5149 VDD.n386 VDD 0.0244044
R5150 VDD.n629 VDD 0.0244044
R5151 VDD.n460 VDD.n459 0.023
R5152 VDD.n499 VDD.n498 0.023
R5153 VDD.n538 VDD.n537 0.023
R5154 VDD.n577 VDD.n576 0.023
R5155 VDD.n985 VDD.n984 0.023
R5156 VDD.n956 VDD.n955 0.023
R5157 VDD.n927 VDD.n926 0.023
R5158 VDD.n898 VDD.n897 0.023
R5159 VDD.n869 VDD.n868 0.023
R5160 VDD.n840 VDD.n839 0.023
R5161 VDD.n128 VDD.n127 0.0222799
R5162 VDD.n143 VDD.n142 0.0222799
R5163 VDD VDD.n0 0.0219868
R5164 VDD.n616 VDD 0.02
R5165 VDD.n465 VDD.n464 0.019
R5166 VDD.n504 VDD.n503 0.019
R5167 VDD.n543 VDD.n542 0.019
R5168 VDD.n582 VDD.n581 0.019
R5169 VDD.n980 VDD.n647 0.019
R5170 VDD.n951 VDD.n675 0.019
R5171 VDD.n922 VDD.n703 0.019
R5172 VDD.n893 VDD.n731 0.019
R5173 VDD.n864 VDD.n759 0.019
R5174 VDD.n835 VDD.n787 0.019
R5175 VDD.n622 VDD.n621 0.0189263
R5176 VDD.n617 VDD.n616 0.0184283
R5177 VDD.n180 VDD.n93 0.0180648
R5178 VDD.n189 VDD.n186 0.0180648
R5179 VDD.n245 VDD.n63 0.0180648
R5180 VDD.n279 VDD.n278 0.0180648
R5181 VDD.n297 VDD.n16 0.0180648
R5182 VDD.n145 VDD 0.0161813
R5183 VDD.n163 VDD.n108 0.014911
R5184 VDD.n193 VDD.n192 0.014911
R5185 VDD.n223 VDD.n73 0.014911
R5186 VDD.n244 VDD.n243 0.014911
R5187 VDD.n296 VDD.n28 0.014911
R5188 VDD.n315 VDD.n314 0.014911
R5189 VDD.n459 VDD.n458 0.0145
R5190 VDD.n498 VDD.n497 0.0145
R5191 VDD.n537 VDD.n536 0.0145
R5192 VDD.n576 VDD.n575 0.0145
R5193 VDD.n615 VDD.n614 0.0145
R5194 VDD.n985 VDD.n645 0.0145
R5195 VDD.n956 VDD.n673 0.0145
R5196 VDD.n927 VDD.n701 0.0145
R5197 VDD.n898 VDD.n729 0.0145
R5198 VDD.n869 VDD.n757 0.0145
R5199 VDD.n840 VDD.n785 0.0145
R5200 VDD.n478 VDD 0.012
R5201 VDD.n517 VDD 0.012
R5202 VDD.n556 VDD 0.012
R5203 VDD.n595 VDD 0.012
R5204 VDD.n632 VDD 0.012
R5205 VDD.n660 VDD 0.012
R5206 VDD.n688 VDD 0.012
R5207 VDD.n716 VDD 0.012
R5208 VDD.n744 VDD 0.012
R5209 VDD.n772 VDD 0.012
R5210 VDD.n800 VDD 0.012
R5211 VDD.n458 VDD 0.0105
R5212 VDD.n497 VDD 0.0105
R5213 VDD.n536 VDD 0.0105
R5214 VDD.n575 VDD 0.0105
R5215 VDD.n614 VDD 0.0105
R5216 VDD.n645 VDD 0.0105
R5217 VDD.n673 VDD 0.0105
R5218 VDD.n701 VDD 0.0105
R5219 VDD.n729 VDD 0.0105
R5220 VDD.n757 VDD 0.0105
R5221 VDD.n785 VDD 0.0105
R5222 VDD VDD.n814 0.01
R5223 VDD VDD.n472 0.009
R5224 VDD.n478 VDD 0.009
R5225 VDD.n477 VDD 0.009
R5226 VDD VDD.n448 0.009
R5227 VDD.n481 VDD 0.009
R5228 VDD VDD.n489 0.009
R5229 VDD VDD.n490 0.009
R5230 VDD.n491 VDD 0.009
R5231 VDD VDD.n511 0.009
R5232 VDD.n517 VDD 0.009
R5233 VDD.n516 VDD 0.009
R5234 VDD VDD.n430 0.009
R5235 VDD.n520 VDD 0.009
R5236 VDD VDD.n528 0.009
R5237 VDD VDD.n529 0.009
R5238 VDD.n530 VDD 0.009
R5239 VDD VDD.n550 0.009
R5240 VDD.n556 VDD 0.009
R5241 VDD.n555 VDD 0.009
R5242 VDD VDD.n412 0.009
R5243 VDD.n559 VDD 0.009
R5244 VDD VDD.n567 0.009
R5245 VDD VDD.n568 0.009
R5246 VDD.n569 VDD 0.009
R5247 VDD VDD.n589 0.009
R5248 VDD.n595 VDD 0.009
R5249 VDD.n594 VDD 0.009
R5250 VDD VDD.n394 0.009
R5251 VDD.n598 VDD 0.009
R5252 VDD VDD.n606 0.009
R5253 VDD VDD.n607 0.009
R5254 VDD.n608 VDD 0.009
R5255 VDD.n632 VDD 0.009
R5256 VDD.n1002 VDD 0.009
R5257 VDD VDD.n1001 0.009
R5258 VDD.n998 VDD 0.009
R5259 VDD.n993 VDD 0.009
R5260 VDD.n992 VDD 0.009
R5261 VDD.n989 VDD 0.009
R5262 VDD.n976 VDD 0.009
R5263 VDD.n660 VDD 0.009
R5264 VDD.n973 VDD 0.009
R5265 VDD VDD.n972 0.009
R5266 VDD.n969 VDD 0.009
R5267 VDD.n964 VDD 0.009
R5268 VDD.n963 VDD 0.009
R5269 VDD.n960 VDD 0.009
R5270 VDD.n947 VDD 0.009
R5271 VDD.n688 VDD 0.009
R5272 VDD.n944 VDD 0.009
R5273 VDD VDD.n943 0.009
R5274 VDD.n940 VDD 0.009
R5275 VDD.n935 VDD 0.009
R5276 VDD.n934 VDD 0.009
R5277 VDD.n931 VDD 0.009
R5278 VDD.n918 VDD 0.009
R5279 VDD.n716 VDD 0.009
R5280 VDD.n915 VDD 0.009
R5281 VDD VDD.n914 0.009
R5282 VDD.n911 VDD 0.009
R5283 VDD.n906 VDD 0.009
R5284 VDD.n905 VDD 0.009
R5285 VDD.n902 VDD 0.009
R5286 VDD.n889 VDD 0.009
R5287 VDD.n744 VDD 0.009
R5288 VDD.n886 VDD 0.009
R5289 VDD VDD.n885 0.009
R5290 VDD.n882 VDD 0.009
R5291 VDD.n877 VDD 0.009
R5292 VDD.n876 VDD 0.009
R5293 VDD.n873 VDD 0.009
R5294 VDD.n860 VDD 0.009
R5295 VDD.n772 VDD 0.009
R5296 VDD.n857 VDD 0.009
R5297 VDD VDD.n856 0.009
R5298 VDD.n853 VDD 0.009
R5299 VDD.n848 VDD 0.009
R5300 VDD.n847 VDD 0.009
R5301 VDD.n844 VDD 0.009
R5302 VDD.n831 VDD 0.009
R5303 VDD.n800 VDD 0.009
R5304 VDD.n828 VDD 0.009
R5305 VDD VDD.n827 0.009
R5306 VDD.n824 VDD 0.009
R5307 VDD.n819 VDD 0.009
R5308 VDD.n818 VDD 0.009
R5309 VDD.n815 VDD 0.009
R5310 VDD VDD.n629 0.00896613
R5311 VDD.n480 VDD.n448 0.0085
R5312 VDD.n519 VDD.n430 0.0085
R5313 VDD.n558 VDD.n412 0.0085
R5314 VDD.n597 VDD.n394 0.0085
R5315 VDD.n1001 VDD.n634 0.0085
R5316 VDD.n972 VDD.n662 0.0085
R5317 VDD.n943 VDD.n690 0.0085
R5318 VDD.n914 VDD.n718 0.0085
R5319 VDD.n885 VDD.n746 0.0085
R5320 VDD.n856 VDD.n774 0.0085
R5321 VDD.n827 VDD.n802 0.0085
R5322 VDD.n490 VDD 0.0075
R5323 VDD.n529 VDD 0.0075
R5324 VDD.n568 VDD 0.0075
R5325 VDD.n607 VDD 0.0075
R5326 VDD VDD.n992 0.0075
R5327 VDD VDD.n963 0.0075
R5328 VDD VDD.n934 0.0075
R5329 VDD VDD.n905 0.0075
R5330 VDD VDD.n876 0.0075
R5331 VDD VDD.n847 0.0075
R5332 VDD VDD.n818 0.0075
R5333 VDD.n814 VDD 0.0065
R5334 VDD.n464 VDD 0.006
R5335 VDD.n503 VDD 0.006
R5336 VDD.n542 VDD 0.006
R5337 VDD.n581 VDD 0.006
R5338 VDD.n980 VDD 0.006
R5339 VDD.n951 VDD 0.006
R5340 VDD.n922 VDD 0.006
R5341 VDD.n893 VDD 0.006
R5342 VDD.n864 VDD 0.006
R5343 VDD.n835 VDD 0.006
R5344 VDD.n621 VDD 0.00597809
R5345 VDD.n475 VDD.n474 0.0055
R5346 VDD.n486 VDD 0.0055
R5347 VDD.n514 VDD.n513 0.0055
R5348 VDD.n525 VDD 0.0055
R5349 VDD.n553 VDD.n552 0.0055
R5350 VDD.n564 VDD 0.0055
R5351 VDD.n592 VDD.n591 0.0055
R5352 VDD.n603 VDD 0.0055
R5353 VDD.n1004 VDD.n630 0.0055
R5354 VDD VDD.n639 0.0055
R5355 VDD.n975 VDD.n658 0.0055
R5356 VDD VDD.n667 0.0055
R5357 VDD.n946 VDD.n686 0.0055
R5358 VDD VDD.n695 0.0055
R5359 VDD.n917 VDD.n714 0.0055
R5360 VDD VDD.n723 0.0055
R5361 VDD.n888 VDD.n742 0.0055
R5362 VDD VDD.n751 0.0055
R5363 VDD.n859 VDD.n770 0.0055
R5364 VDD VDD.n779 0.0055
R5365 VDD.n830 VDD.n798 0.0055
R5366 VDD VDD.n807 0.0055
R5367 VDD.n616 VDD.n615 0.005
R5368 VDD.n474 VDD 0.004
R5369 VDD.n487 VDD.n486 0.004
R5370 VDD.n513 VDD 0.004
R5371 VDD.n526 VDD.n525 0.004
R5372 VDD.n552 VDD 0.004
R5373 VDD.n565 VDD.n564 0.004
R5374 VDD.n591 VDD 0.004
R5375 VDD.n604 VDD.n603 0.004
R5376 VDD VDD.n630 0.004
R5377 VDD.n997 VDD.n639 0.004
R5378 VDD VDD.n658 0.004
R5379 VDD.n968 VDD.n667 0.004
R5380 VDD VDD.n686 0.004
R5381 VDD.n939 VDD.n695 0.004
R5382 VDD VDD.n714 0.004
R5383 VDD.n910 VDD.n723 0.004
R5384 VDD VDD.n742 0.004
R5385 VDD.n881 VDD.n751 0.004
R5386 VDD VDD.n770 0.004
R5387 VDD.n852 VDD.n779 0.004
R5388 VDD VDD.n798 0.004
R5389 VDD.n823 VDD.n807 0.004
R5390 VDD VDD.n477 0.003
R5391 VDD VDD.n516 0.003
R5392 VDD VDD.n555 0.003
R5393 VDD VDD.n594 0.003
R5394 VDD.n1002 VDD 0.003
R5395 VDD.n973 VDD 0.003
R5396 VDD.n944 VDD 0.003
R5397 VDD.n915 VDD 0.003
R5398 VDD.n886 VDD 0.003
R5399 VDD.n857 VDD 0.003
R5400 VDD.n828 VDD 0.003
R5401 VDD.n460 VDD 0.002
R5402 VDD.n499 VDD 0.002
R5403 VDD.n538 VDD 0.002
R5404 VDD.n577 VDD 0.002
R5405 VDD.n984 VDD 0.002
R5406 VDD.n955 VDD 0.002
R5407 VDD.n926 VDD 0.002
R5408 VDD.n897 VDD 0.002
R5409 VDD.n868 VDD 0.002
R5410 VDD.n839 VDD 0.002
R5411 VDD.n617 VDD 0.00199402
R5412 VDD VDD.n480 0.001
R5413 VDD VDD.n519 0.001
R5414 VDD VDD.n558 0.001
R5415 VDD VDD.n597 0.001
R5416 VDD VDD.n634 0.001
R5417 VDD VDD.n662 0.001
R5418 VDD VDD.n690 0.001
R5419 VDD VDD.n718 0.001
R5420 VDD VDD.n746 0.001
R5421 VDD VDD.n774 0.001
R5422 VDD VDD.n802 0.001
R5423 ia_opamp_0.V2.n35 ia_opamp_0.V2.t38 492.029
R5424 ia_opamp_0.V2.n38 ia_opamp_0.V2.t12 39.1599
R5425 ia_opamp_0.V2.n0 ia_opamp_0.V2.t13 21.5504
R5426 ia_opamp_0.V2.n1 ia_opamp_0.V2.t0 21.4819
R5427 ia_opamp_0.V2.n0 ia_opamp_0.V2.t6 21.4809
R5428 ia_opamp_0.V2.n2 ia_opamp_0.V2.t32 21.4809
R5429 ia_opamp_0.V2.n3 ia_opamp_0.V2.t21 21.4809
R5430 ia_opamp_0.V2.n4 ia_opamp_0.V2.t23 21.4809
R5431 ia_opamp_0.V2.n5 ia_opamp_0.V2.t2 21.4809
R5432 ia_opamp_0.V2.n6 ia_opamp_0.V2.t14 21.4809
R5433 ia_opamp_0.V2.n7 ia_opamp_0.V2.t29 21.4809
R5434 ia_opamp_0.V2.n8 ia_opamp_0.V2.t1 21.4809
R5435 ia_opamp_0.V2.n9 ia_opamp_0.V2.t3 21.4809
R5436 ia_opamp_0.V2.n10 ia_opamp_0.V2.t7 21.4809
R5437 ia_opamp_0.V2.n11 ia_opamp_0.V2.t22 21.4809
R5438 ia_opamp_0.V2.n12 ia_opamp_0.V2.t4 21.4809
R5439 ia_opamp_0.V2.n13 ia_opamp_0.V2.t8 21.4809
R5440 ia_opamp_0.V2.n14 ia_opamp_0.V2.t17 21.4809
R5441 ia_opamp_0.V2.n15 ia_opamp_0.V2.t30 21.4809
R5442 ia_opamp_0.V2.n16 ia_opamp_0.V2.t16 21.4809
R5443 ia_opamp_0.V2.n17 ia_opamp_0.V2.t19 21.4809
R5444 ia_opamp_0.V2.n18 ia_opamp_0.V2.t27 21.4809
R5445 ia_opamp_0.V2.n19 ia_opamp_0.V2.t18 21.4809
R5446 ia_opamp_0.V2.n20 ia_opamp_0.V2.t24 21.4809
R5447 ia_opamp_0.V2.n21 ia_opamp_0.V2.t20 21.4809
R5448 ia_opamp_0.V2.n22 ia_opamp_0.V2.t10 21.4809
R5449 ia_opamp_0.V2.n23 ia_opamp_0.V2.t9 21.4809
R5450 ia_opamp_0.V2.n24 ia_opamp_0.V2.t5 21.4809
R5451 ia_opamp_0.V2.n25 ia_opamp_0.V2.t31 21.4809
R5452 ia_opamp_0.V2.n26 ia_opamp_0.V2.t26 21.4809
R5453 ia_opamp_0.V2.n27 ia_opamp_0.V2.t15 21.4809
R5454 ia_opamp_0.V2.n28 ia_opamp_0.V2.t25 21.4809
R5455 ia_opamp_0.V2.n29 ia_opamp_0.V2.t28 21.4809
R5456 ia_opamp_0.V2.n30 ia_opamp_0.V2.t33 21.4809
R5457 ia_opamp_0.V2.n33 ia_opamp_0.V2.n31 13.4669
R5458 ia_opamp_0.V2.n33 ia_opamp_0.V2.n32 13.3799
R5459 ia_opamp_0.V2.n40 ia_opamp_0.V2.n39 8.26762
R5460 ia_opamp_0.V2.n37 ia_opamp_0.V2.n36 6.92437
R5461 ia_opamp_0.V2.n39 ia_opamp_0.V2.n38 5.93365
R5462 ia_opamp_0.V2.n38 ia_opamp_0.V2.t11 4.35292
R5463 ia_opamp_0.V2.n34 ia_opamp_0.V2 2.58592
R5464 ia_opamp_0.V2.n34 ia_opamp_0.V2.n33 2.00817
R5465 ia_opamp_0.V2.n31 ia_opamp_0.V2.t35 1.45813
R5466 ia_opamp_0.V2.n31 ia_opamp_0.V2.t36 1.45813
R5467 ia_opamp_0.V2.n32 ia_opamp_0.V2.t34 1.45813
R5468 ia_opamp_0.V2.n32 ia_opamp_0.V2.t37 1.45813
R5469 ia_opamp_0.V2 ia_opamp_0.V2.n40 0.419948
R5470 ia_opamp_0.V2.n37 ia_opamp_0.V2.n34 0.227129
R5471 ia_opamp_0.V2.n23 ia_opamp_0.V2.n22 0.223778
R5472 ia_opamp_0.V2.n27 ia_opamp_0.V2.n26 0.205963
R5473 ia_opamp_0.V2.n15 ia_opamp_0.V2.n14 0.196462
R5474 ia_opamp_0.V2.n29 ia_opamp_0.V2.n28 0.188148
R5475 ia_opamp_0.V2.n39 ia_opamp_0.V2.n37 0.167924
R5476 ia_opamp_0.V2.n30 ia_opamp_0.V2.n29 0.15727
R5477 ia_opamp_0.V2.n35 ia_opamp_0.V2 0.0796667
R5478 ia_opamp_0.V2.n1 ia_opamp_0.V2.n0 0.0699774
R5479 ia_opamp_0.V2.n2 ia_opamp_0.V2.n1 0.0699774
R5480 ia_opamp_0.V2.n3 ia_opamp_0.V2.n2 0.0699774
R5481 ia_opamp_0.V2.n4 ia_opamp_0.V2.n3 0.0699774
R5482 ia_opamp_0.V2.n5 ia_opamp_0.V2.n4 0.0699774
R5483 ia_opamp_0.V2.n6 ia_opamp_0.V2.n5 0.0699774
R5484 ia_opamp_0.V2.n7 ia_opamp_0.V2.n6 0.0699774
R5485 ia_opamp_0.V2.n8 ia_opamp_0.V2.n7 0.0699774
R5486 ia_opamp_0.V2.n9 ia_opamp_0.V2.n8 0.0699774
R5487 ia_opamp_0.V2.n10 ia_opamp_0.V2.n9 0.0699774
R5488 ia_opamp_0.V2.n11 ia_opamp_0.V2.n10 0.0699774
R5489 ia_opamp_0.V2.n12 ia_opamp_0.V2.n11 0.0699774
R5490 ia_opamp_0.V2.n13 ia_opamp_0.V2.n12 0.0699774
R5491 ia_opamp_0.V2.n14 ia_opamp_0.V2.n13 0.0699774
R5492 ia_opamp_0.V2.n16 ia_opamp_0.V2.n15 0.0699774
R5493 ia_opamp_0.V2.n17 ia_opamp_0.V2.n16 0.0699774
R5494 ia_opamp_0.V2.n18 ia_opamp_0.V2.n17 0.0699774
R5495 ia_opamp_0.V2.n19 ia_opamp_0.V2.n18 0.0699774
R5496 ia_opamp_0.V2.n20 ia_opamp_0.V2.n19 0.0699774
R5497 ia_opamp_0.V2.n21 ia_opamp_0.V2.n20 0.0699774
R5498 ia_opamp_0.V2.n22 ia_opamp_0.V2.n21 0.0699774
R5499 ia_opamp_0.V2.n24 ia_opamp_0.V2.n23 0.0699774
R5500 ia_opamp_0.V2.n25 ia_opamp_0.V2.n24 0.0699774
R5501 ia_opamp_0.V2.n26 ia_opamp_0.V2.n25 0.0699774
R5502 ia_opamp_0.V2.n28 ia_opamp_0.V2.n27 0.0699774
R5503 ia_opamp_0.V2.n36 ia_opamp_0.V2.n35 0.0686818
R5504 ia_opamp_0.V2.n36 ia_opamp_0.V2 0.0108306
R5505 ia_opamp_0.V2.n40 ia_opamp_0.V2.n30 0.000796912
R5506 DVSS.n2784 DVSS.t2 20051.8
R5507 DVSS.n1722 DVSS.n518 5082
R5508 DVSS.n696 DVSS.n578 5082
R5509 DVSS.n1341 DVSS.n1340 5082
R5510 DVSS.n1170 DVSS.n1169 5082
R5511 DVSS.n988 DVSS.n987 5082
R5512 DVSS.n1840 DVSS.n1839 5082
R5513 DVSS.n2022 DVSS.n2021 5082
R5514 DVSS.n2204 DVSS.n2203 5082
R5515 DVSS.n2375 DVSS.n2374 5082
R5516 DVSS.n204 DVSS.n86 5082
R5517 DVSS.n2715 DVSS.n26 5082
R5518 DVSS.n1754 DVSS.t176 5042.05
R5519 DVSS.n1653 DVSS.t229 5042.05
R5520 DVSS.n671 DVSS.t146 5042.05
R5521 DVSS.n1261 DVSS.t196 5042.05
R5522 DVSS.n1079 DVSS.t170 5042.05
R5523 DVSS.n1931 DVSS.t237 5042.05
R5524 DVSS.n2113 DVSS.t182 5042.05
R5525 DVSS.n2295 DVSS.t138 5042.05
R5526 DVSS.n179 DVSS.t126 5042.05
R5527 DVSS.n2646 DVSS.t88 5042.05
R5528 DVSS.n2747 DVSS.t22 5042.05
R5529 DVSS.n2785 DVSS.n2784 1739.72
R5530 DVSS.n904 DVSS.t269 1435.41
R5531 DVSS.n954 DVSS.n953 1118.03
R5532 DVSS.n1077 DVSS.n1076 979.885
R5533 DVSS.n1259 DVSS.n1258 979.885
R5534 DVSS.n1427 DVSS.n1426 979.885
R5535 DVSS.n1651 DVSS.n546 979.885
R5536 DVSS.n1590 DVSS.n1584 979.885
R5537 DVSS.n1929 DVSS.n1928 979.885
R5538 DVSS.n2111 DVSS.n2110 979.885
R5539 DVSS.n2293 DVSS.n2292 979.885
R5540 DVSS.n2461 DVSS.n2460 979.885
R5541 DVSS.n2644 DVSS.n54 979.885
R5542 DVSS.n989 DVSS.n896 898.723
R5543 DVSS.n998 DVSS.n891 898.723
R5544 DVSS.n999 DVSS.n998 898.723
R5545 DVSS.n1171 DVSS.n824 898.723
R5546 DVSS.n1180 DVSS.n819 898.723
R5547 DVSS.n1181 DVSS.n1180 898.723
R5548 DVSS.n1342 DVSS.n623 898.723
R5549 DVSS.n1351 DVSS.n618 898.723
R5550 DVSS.n1352 DVSS.n1351 898.723
R5551 DVSS.n1429 DVSS.n1428 898.723
R5552 DVSS.n1439 DVSS.n1438 898.723
R5553 DVSS.n1441 DVSS.n1439 898.723
R5554 DVSS.n1650 DVSS.n547 898.723
R5555 DVSS.n1567 DVSS.n1566 898.723
R5556 DVSS.n1569 DVSS.n1567 898.723
R5557 DVSS.n1841 DVSS.n476 898.723
R5558 DVSS.n1850 DVSS.n471 898.723
R5559 DVSS.n1851 DVSS.n1850 898.723
R5560 DVSS.n2023 DVSS.n404 898.723
R5561 DVSS.n2032 DVSS.n399 898.723
R5562 DVSS.n2033 DVSS.n2032 898.723
R5563 DVSS.n2205 DVSS.n332 898.723
R5564 DVSS.n2214 DVSS.n327 898.723
R5565 DVSS.n2215 DVSS.n2214 898.723
R5566 DVSS.n2376 DVSS.n131 898.723
R5567 DVSS.n2385 DVSS.n126 898.723
R5568 DVSS.n2386 DVSS.n2385 898.723
R5569 DVSS.n2463 DVSS.n2462 898.723
R5570 DVSS.n2473 DVSS.n2472 898.723
R5571 DVSS.n2475 DVSS.n2473 898.723
R5572 DVSS.n2643 DVSS.n55 898.723
R5573 DVSS.n2564 DVSS.n2563 898.723
R5574 DVSS.n2566 DVSS.n2564 898.723
R5575 DVSS.n2763 DVSS.n5 769.572
R5576 DVSS.n916 DVSS.n914 769.572
R5577 DVSS.n2786 DVSS.n2785 769.572
R5578 DVSS.n932 DVSS.n905 769.572
R5579 DVSS.n954 DVSS.n896 748.937
R5580 DVSS.n1077 DVSS.n824 748.937
R5581 DVSS.n1259 DVSS.n623 748.937
R5582 DVSS.n1429 DVSS.n1427 748.937
R5583 DVSS.n1651 DVSS.n1650 748.937
R5584 DVSS.n1584 DVSS.n476 748.937
R5585 DVSS.n1929 DVSS.n404 748.937
R5586 DVSS.n2111 DVSS.n332 748.937
R5587 DVSS.n2293 DVSS.n131 748.937
R5588 DVSS.n2463 DVSS.n2461 748.937
R5589 DVSS.n2644 DVSS.n2643 748.937
R5590 DVSS.t2 DVSS.n2783 704.931
R5591 DVSS.n988 DVSS.n891 674.043
R5592 DVSS.n1170 DVSS.n819 674.043
R5593 DVSS.n1341 DVSS.n618 674.043
R5594 DVSS.n1438 DVSS.n578 674.043
R5595 DVSS.n1566 DVSS.n518 674.043
R5596 DVSS.n1840 DVSS.n471 674.043
R5597 DVSS.n2022 DVSS.n399 674.043
R5598 DVSS.n2204 DVSS.n327 674.043
R5599 DVSS.n2375 DVSS.n126 674.043
R5600 DVSS.n2472 DVSS.n86 674.043
R5601 DVSS.n2563 DVSS.n26 674.043
R5602 DVSS.n1077 DVSS.n858 623.971
R5603 DVSS.n1259 DVSS.n786 623.971
R5604 DVSS.n1427 DVSS.n584 623.971
R5605 DVSS.n1651 DVSS.n545 623.971
R5606 DVSS.n1584 DVSS.n1583 623.971
R5607 DVSS.n1929 DVSS.n438 623.971
R5608 DVSS.n2111 DVSS.n366 623.971
R5609 DVSS.n2293 DVSS.n294 623.971
R5610 DVSS.n2461 DVSS.n92 623.971
R5611 DVSS.n2644 DVSS.n53 623.971
R5612 DVSS.n2784 DVSS.n3 623.971
R5613 DVSS.n2760 DVSS.n2759 585
R5614 DVSS.n2771 DVSS.n2758 585
R5615 DVSS.n2772 DVSS.n2757 585
R5616 DVSS.n2756 DVSS.n2755 585
R5617 DVSS.n2776 DVSS.n2754 585
R5618 DVSS.n2777 DVSS.n2753 585
R5619 DVSS.n12 DVSS.n10 585
R5620 DVSS.n2782 DVSS.n2781 585
R5621 DVSS.n2783 DVSS.n2782 585
R5622 DVSS.n11 DVSS.n9 585
R5623 DVSS.n9 DVSS.n4 585
R5624 DVSS.n2750 DVSS.n2749 585
R5625 DVSS.n2749 DVSS.n2748 585
R5626 DVSS.n14 DVSS.n13 585
R5627 DVSS.n2746 DVSS.n14 585
R5628 DVSS.n2744 DVSS.n2743 585
R5629 DVSS.n2745 DVSS.n2744 585
R5630 DVSS.n17 DVSS.n16 585
R5631 DVSS.n16 DVSS.n15 585
R5632 DVSS.n2726 DVSS.n2721 585
R5633 DVSS.n2721 DVSS.n2720 585
R5634 DVSS.n2727 DVSS.n25 585
R5635 DVSS.n2719 DVSS.n25 585
R5636 DVSS.n2717 DVSS.n24 585
R5637 DVSS.n2718 DVSS.n2717 585
R5638 DVSS.n2731 DVSS.n23 585
R5639 DVSS.n2716 DVSS.n23 585
R5640 DVSS.n2732 DVSS.n22 585
R5641 DVSS.n2714 DVSS.n22 585
R5642 DVSS.n2712 DVSS.n21 585
R5643 DVSS.n2713 DVSS.n2712 585
R5644 DVSS.n2711 DVSS.n2710 585
R5645 DVSS.n2711 DVSS.n27 585
R5646 DVSS.n29 DVSS.n28 585
R5647 DVSS.n2702 DVSS.n28 585
R5648 DVSS.n2705 DVSS.n2704 585
R5649 DVSS.n2704 DVSS.n2703 585
R5650 DVSS.n31 DVSS.n30 585
R5651 DVSS.n2701 DVSS.n31 585
R5652 DVSS.n2699 DVSS.n2698 585
R5653 DVSS.n2700 DVSS.n2699 585
R5654 DVSS.n34 DVSS.n33 585
R5655 DVSS.n33 DVSS.n32 585
R5656 DVSS.n2693 DVSS.n2692 585
R5657 DVSS.n2692 DVSS.n2691 585
R5658 DVSS.n36 DVSS.n35 585
R5659 DVSS.n2690 DVSS.n36 585
R5660 DVSS.n2688 DVSS.n2687 585
R5661 DVSS.n2689 DVSS.n2688 585
R5662 DVSS.n38 DVSS.n37 585
R5663 DVSS.n2674 DVSS.n37 585
R5664 DVSS.n2677 DVSS.n2676 585
R5665 DVSS.n2676 DVSS.n2675 585
R5666 DVSS.n40 DVSS.n39 585
R5667 DVSS.n2673 DVSS.n40 585
R5668 DVSS.n2671 DVSS.n2670 585
R5669 DVSS.n2672 DVSS.n2671 585
R5670 DVSS.n43 DVSS.n42 585
R5671 DVSS.n42 DVSS.n41 585
R5672 DVSS.n2665 DVSS.n2664 585
R5673 DVSS.n2664 DVSS.n2663 585
R5674 DVSS.n45 DVSS.n44 585
R5675 DVSS.n2662 DVSS.n45 585
R5676 DVSS.n2660 DVSS.n2659 585
R5677 DVSS.n2661 DVSS.n2660 585
R5678 DVSS.n47 DVSS.n46 585
R5679 DVSS.n2647 DVSS.n46 585
R5680 DVSS.n2650 DVSS.n2649 585
R5681 DVSS.n2649 DVSS.n2648 585
R5682 DVSS.n50 DVSS.n49 585
R5683 DVSS.n51 DVSS.n50 585
R5684 DVSS.n211 DVSS.n210 585
R5685 DVSS.n210 DVSS.n209 585
R5686 DVSS.n219 DVSS.n166 585
R5687 DVSS.n208 DVSS.n166 585
R5688 DVSS.n220 DVSS.n165 585
R5689 DVSS.n207 DVSS.n165 585
R5690 DVSS.n205 DVSS.n164 585
R5691 DVSS.n206 DVSS.n205 585
R5692 DVSS.n227 DVSS.n163 585
R5693 DVSS.n203 DVSS.n163 585
R5694 DVSS.n228 DVSS.n162 585
R5695 DVSS.n202 DVSS.n162 585
R5696 DVSS.n200 DVSS.n161 585
R5697 DVSS.n201 DVSS.n200 585
R5698 DVSS.n232 DVSS.n160 585
R5699 DVSS.n199 DVSS.n160 585
R5700 DVSS.n233 DVSS.n159 585
R5701 DVSS.n198 DVSS.n159 585
R5702 DVSS.n196 DVSS.n158 585
R5703 DVSS.n197 DVSS.n196 585
R5704 DVSS.n237 DVSS.n157 585
R5705 DVSS.n195 DVSS.n157 585
R5706 DVSS.n238 DVSS.n156 585
R5707 DVSS.n194 DVSS.n156 585
R5708 DVSS.n241 DVSS.n155 585
R5709 DVSS.n193 DVSS.n155 585
R5710 DVSS.n242 DVSS.n154 585
R5711 DVSS.n192 DVSS.n154 585
R5712 DVSS.n190 DVSS.n152 585
R5713 DVSS.n191 DVSS.n190 585
R5714 DVSS.n250 DVSS.n151 585
R5715 DVSS.n189 DVSS.n151 585
R5716 DVSS.n251 DVSS.n150 585
R5717 DVSS.n188 DVSS.n150 585
R5718 DVSS.n186 DVSS.n149 585
R5719 DVSS.n187 DVSS.n186 585
R5720 DVSS.n255 DVSS.n148 585
R5721 DVSS.n185 DVSS.n148 585
R5722 DVSS.n256 DVSS.n147 585
R5723 DVSS.n184 DVSS.n147 585
R5724 DVSS.n182 DVSS.n146 585
R5725 DVSS.n183 DVSS.n182 585
R5726 DVSS.n260 DVSS.n145 585
R5727 DVSS.n181 DVSS.n145 585
R5728 DVSS.n261 DVSS.n144 585
R5729 DVSS.n180 DVSS.n144 585
R5730 DVSS.n177 DVSS.n143 585
R5731 DVSS.n178 DVSS.n177 585
R5732 DVSS.n176 DVSS.n170 585
R5733 DVSS.n176 DVSS.n175 585
R5734 DVSS.n167 DVSS.n139 585
R5735 DVSS.n174 DVSS.n167 585
R5736 DVSS.n2366 DVSS.n138 585
R5737 DVSS.n173 DVSS.n138 585
R5738 DVSS.n2367 DVSS.n137 585
R5739 DVSS.n172 DVSS.n137 585
R5740 DVSS.n136 DVSS.n134 585
R5741 DVSS.n171 DVSS.n134 585
R5742 DVSS.n2372 DVSS.n2371 585
R5743 DVSS.n2373 DVSS.n2372 585
R5744 DVSS.n135 DVSS.n133 585
R5745 DVSS.n133 DVSS.n132 585
R5746 DVSS.n2355 DVSS.n2354 585
R5747 DVSS.n2354 DVSS.n2353 585
R5748 DVSS.n267 DVSS.n266 585
R5749 DVSS.n2352 DVSS.n267 585
R5750 DVSS.n2350 DVSS.n2349 585
R5751 DVSS.n2351 DVSS.n2350 585
R5752 DVSS.n270 DVSS.n269 585
R5753 DVSS.n269 DVSS.n268 585
R5754 DVSS.n2344 DVSS.n2343 585
R5755 DVSS.n2343 DVSS.n2342 585
R5756 DVSS.n272 DVSS.n271 585
R5757 DVSS.n2341 DVSS.n272 585
R5758 DVSS.n2339 DVSS.n2338 585
R5759 DVSS.n2340 DVSS.n2339 585
R5760 DVSS.n2334 DVSS.n274 585
R5761 DVSS.n274 DVSS.n273 585
R5762 DVSS.n2333 DVSS.n276 585
R5763 DVSS.n2322 DVSS.n276 585
R5764 DVSS.n281 DVSS.n275 585
R5765 DVSS.n2323 DVSS.n281 585
R5766 DVSS.n2326 DVSS.n2325 585
R5767 DVSS.n2325 DVSS.n2324 585
R5768 DVSS.n280 DVSS.n279 585
R5769 DVSS.n2321 DVSS.n280 585
R5770 DVSS.n2319 DVSS.n2318 585
R5771 DVSS.n2320 DVSS.n2319 585
R5772 DVSS.n284 DVSS.n283 585
R5773 DVSS.n283 DVSS.n282 585
R5774 DVSS.n2313 DVSS.n2312 585
R5775 DVSS.n2312 DVSS.n2311 585
R5776 DVSS.n286 DVSS.n285 585
R5777 DVSS.n2310 DVSS.n286 585
R5778 DVSS.n2308 DVSS.n2307 585
R5779 DVSS.n2309 DVSS.n2308 585
R5780 DVSS.n289 DVSS.n288 585
R5781 DVSS.n288 DVSS.n287 585
R5782 DVSS.n2298 DVSS.n2297 585
R5783 DVSS.n2297 DVSS.n2296 585
R5784 DVSS.n292 DVSS.n291 585
R5785 DVSS.n2184 DVSS.n292 585
R5786 DVSS.n2187 DVSS.n2186 585
R5787 DVSS.n2186 DVSS.n2185 585
R5788 DVSS.n2195 DVSS.n2180 585
R5789 DVSS.n2183 DVSS.n2180 585
R5790 DVSS.n2196 DVSS.n2179 585
R5791 DVSS.n2182 DVSS.n2179 585
R5792 DVSS.n337 DVSS.n335 585
R5793 DVSS.n2181 DVSS.n335 585
R5794 DVSS.n2201 DVSS.n2200 585
R5795 DVSS.n2202 DVSS.n2201 585
R5796 DVSS.n336 DVSS.n334 585
R5797 DVSS.n334 DVSS.n333 585
R5798 DVSS.n2173 DVSS.n2172 585
R5799 DVSS.n2172 DVSS.n2171 585
R5800 DVSS.n339 DVSS.n338 585
R5801 DVSS.n2170 DVSS.n339 585
R5802 DVSS.n2168 DVSS.n2167 585
R5803 DVSS.n2169 DVSS.n2168 585
R5804 DVSS.n342 DVSS.n341 585
R5805 DVSS.n341 DVSS.n340 585
R5806 DVSS.n2162 DVSS.n2161 585
R5807 DVSS.n2161 DVSS.n2160 585
R5808 DVSS.n344 DVSS.n343 585
R5809 DVSS.n2159 DVSS.n344 585
R5810 DVSS.n2157 DVSS.n2156 585
R5811 DVSS.n2158 DVSS.n2157 585
R5812 DVSS.n2152 DVSS.n346 585
R5813 DVSS.n346 DVSS.n345 585
R5814 DVSS.n2151 DVSS.n348 585
R5815 DVSS.n2140 DVSS.n348 585
R5816 DVSS.n353 DVSS.n347 585
R5817 DVSS.n2141 DVSS.n353 585
R5818 DVSS.n2144 DVSS.n2143 585
R5819 DVSS.n2143 DVSS.n2142 585
R5820 DVSS.n352 DVSS.n351 585
R5821 DVSS.n2139 DVSS.n352 585
R5822 DVSS.n2137 DVSS.n2136 585
R5823 DVSS.n2138 DVSS.n2137 585
R5824 DVSS.n356 DVSS.n355 585
R5825 DVSS.n355 DVSS.n354 585
R5826 DVSS.n2131 DVSS.n2130 585
R5827 DVSS.n2130 DVSS.n2129 585
R5828 DVSS.n358 DVSS.n357 585
R5829 DVSS.n2128 DVSS.n358 585
R5830 DVSS.n2126 DVSS.n2125 585
R5831 DVSS.n2127 DVSS.n2126 585
R5832 DVSS.n361 DVSS.n360 585
R5833 DVSS.n360 DVSS.n359 585
R5834 DVSS.n2116 DVSS.n2115 585
R5835 DVSS.n2115 DVSS.n2114 585
R5836 DVSS.n364 DVSS.n363 585
R5837 DVSS.n2002 DVSS.n364 585
R5838 DVSS.n2005 DVSS.n2004 585
R5839 DVSS.n2004 DVSS.n2003 585
R5840 DVSS.n2013 DVSS.n1998 585
R5841 DVSS.n2001 DVSS.n1998 585
R5842 DVSS.n2014 DVSS.n1997 585
R5843 DVSS.n2000 DVSS.n1997 585
R5844 DVSS.n409 DVSS.n407 585
R5845 DVSS.n1999 DVSS.n407 585
R5846 DVSS.n2019 DVSS.n2018 585
R5847 DVSS.n2020 DVSS.n2019 585
R5848 DVSS.n408 DVSS.n406 585
R5849 DVSS.n406 DVSS.n405 585
R5850 DVSS.n1991 DVSS.n1990 585
R5851 DVSS.n1990 DVSS.n1989 585
R5852 DVSS.n411 DVSS.n410 585
R5853 DVSS.n1988 DVSS.n411 585
R5854 DVSS.n1986 DVSS.n1985 585
R5855 DVSS.n1987 DVSS.n1986 585
R5856 DVSS.n414 DVSS.n413 585
R5857 DVSS.n413 DVSS.n412 585
R5858 DVSS.n1980 DVSS.n1979 585
R5859 DVSS.n1979 DVSS.n1978 585
R5860 DVSS.n416 DVSS.n415 585
R5861 DVSS.n1977 DVSS.n416 585
R5862 DVSS.n1975 DVSS.n1974 585
R5863 DVSS.n1976 DVSS.n1975 585
R5864 DVSS.n1970 DVSS.n418 585
R5865 DVSS.n418 DVSS.n417 585
R5866 DVSS.n1969 DVSS.n420 585
R5867 DVSS.n1958 DVSS.n420 585
R5868 DVSS.n425 DVSS.n419 585
R5869 DVSS.n1959 DVSS.n425 585
R5870 DVSS.n1962 DVSS.n1961 585
R5871 DVSS.n1961 DVSS.n1960 585
R5872 DVSS.n424 DVSS.n423 585
R5873 DVSS.n1957 DVSS.n424 585
R5874 DVSS.n1955 DVSS.n1954 585
R5875 DVSS.n1956 DVSS.n1955 585
R5876 DVSS.n428 DVSS.n427 585
R5877 DVSS.n427 DVSS.n426 585
R5878 DVSS.n1949 DVSS.n1948 585
R5879 DVSS.n1948 DVSS.n1947 585
R5880 DVSS.n430 DVSS.n429 585
R5881 DVSS.n1946 DVSS.n430 585
R5882 DVSS.n1944 DVSS.n1943 585
R5883 DVSS.n1945 DVSS.n1944 585
R5884 DVSS.n433 DVSS.n432 585
R5885 DVSS.n432 DVSS.n431 585
R5886 DVSS.n1934 DVSS.n1933 585
R5887 DVSS.n1933 DVSS.n1932 585
R5888 DVSS.n436 DVSS.n435 585
R5889 DVSS.n1820 DVSS.n436 585
R5890 DVSS.n1823 DVSS.n1822 585
R5891 DVSS.n1822 DVSS.n1821 585
R5892 DVSS.n1831 DVSS.n1816 585
R5893 DVSS.n1819 DVSS.n1816 585
R5894 DVSS.n1832 DVSS.n1815 585
R5895 DVSS.n1818 DVSS.n1815 585
R5896 DVSS.n481 DVSS.n479 585
R5897 DVSS.n1817 DVSS.n479 585
R5898 DVSS.n1837 DVSS.n1836 585
R5899 DVSS.n1838 DVSS.n1837 585
R5900 DVSS.n480 DVSS.n478 585
R5901 DVSS.n478 DVSS.n477 585
R5902 DVSS.n1809 DVSS.n1808 585
R5903 DVSS.n1808 DVSS.n1807 585
R5904 DVSS.n483 DVSS.n482 585
R5905 DVSS.n1806 DVSS.n483 585
R5906 DVSS.n1804 DVSS.n1803 585
R5907 DVSS.n1805 DVSS.n1804 585
R5908 DVSS.n486 DVSS.n485 585
R5909 DVSS.n485 DVSS.n484 585
R5910 DVSS.n1798 DVSS.n1797 585
R5911 DVSS.n1797 DVSS.n1796 585
R5912 DVSS.n488 DVSS.n487 585
R5913 DVSS.n1795 DVSS.n488 585
R5914 DVSS.n1793 DVSS.n1792 585
R5915 DVSS.n1794 DVSS.n1793 585
R5916 DVSS.n1788 DVSS.n490 585
R5917 DVSS.n490 DVSS.n489 585
R5918 DVSS.n1787 DVSS.n492 585
R5919 DVSS.n1777 DVSS.n492 585
R5920 DVSS.n1781 DVSS.n1780 585
R5921 DVSS.n1780 DVSS.n1779 585
R5922 DVSS.n496 DVSS.n495 585
R5923 DVSS.n1776 DVSS.n496 585
R5924 DVSS.n1774 DVSS.n1773 585
R5925 DVSS.n1775 DVSS.n1774 585
R5926 DVSS.n499 DVSS.n498 585
R5927 DVSS.n498 DVSS.n497 585
R5928 DVSS.n1768 DVSS.n1767 585
R5929 DVSS.n1767 DVSS.n1766 585
R5930 DVSS.n501 DVSS.n500 585
R5931 DVSS.n1765 DVSS.n501 585
R5932 DVSS.n1763 DVSS.n1762 585
R5933 DVSS.n1764 DVSS.n1763 585
R5934 DVSS.n504 DVSS.n503 585
R5935 DVSS.n503 DVSS.n502 585
R5936 DVSS.n1757 DVSS.n1756 585
R5937 DVSS.n1756 DVSS.n1755 585
R5938 DVSS.n506 DVSS.n505 585
R5939 DVSS.n1753 DVSS.n506 585
R5940 DVSS.n1751 DVSS.n1750 585
R5941 DVSS.n1752 DVSS.n1751 585
R5942 DVSS.n509 DVSS.n508 585
R5943 DVSS.n508 DVSS.n507 585
R5944 DVSS.n1733 DVSS.n1728 585
R5945 DVSS.n1728 DVSS.n1727 585
R5946 DVSS.n1734 DVSS.n517 585
R5947 DVSS.n1726 DVSS.n517 585
R5948 DVSS.n1724 DVSS.n516 585
R5949 DVSS.n1725 DVSS.n1724 585
R5950 DVSS.n1738 DVSS.n515 585
R5951 DVSS.n1723 DVSS.n515 585
R5952 DVSS.n1739 DVSS.n514 585
R5953 DVSS.n1721 DVSS.n514 585
R5954 DVSS.n1719 DVSS.n513 585
R5955 DVSS.n1720 DVSS.n1719 585
R5956 DVSS.n1718 DVSS.n1717 585
R5957 DVSS.n1718 DVSS.n519 585
R5958 DVSS.n521 DVSS.n520 585
R5959 DVSS.n1709 DVSS.n520 585
R5960 DVSS.n1712 DVSS.n1711 585
R5961 DVSS.n1711 DVSS.n1710 585
R5962 DVSS.n523 DVSS.n522 585
R5963 DVSS.n1708 DVSS.n523 585
R5964 DVSS.n1706 DVSS.n1705 585
R5965 DVSS.n1707 DVSS.n1706 585
R5966 DVSS.n526 DVSS.n525 585
R5967 DVSS.n525 DVSS.n524 585
R5968 DVSS.n1700 DVSS.n1699 585
R5969 DVSS.n1699 DVSS.n1698 585
R5970 DVSS.n528 DVSS.n527 585
R5971 DVSS.n1697 DVSS.n528 585
R5972 DVSS.n1695 DVSS.n1694 585
R5973 DVSS.n1696 DVSS.n1695 585
R5974 DVSS.n530 DVSS.n529 585
R5975 DVSS.n1681 DVSS.n529 585
R5976 DVSS.n1684 DVSS.n1683 585
R5977 DVSS.n1683 DVSS.n1682 585
R5978 DVSS.n532 DVSS.n531 585
R5979 DVSS.n1680 DVSS.n532 585
R5980 DVSS.n1678 DVSS.n1677 585
R5981 DVSS.n1679 DVSS.n1678 585
R5982 DVSS.n535 DVSS.n534 585
R5983 DVSS.n534 DVSS.n533 585
R5984 DVSS.n1672 DVSS.n1671 585
R5985 DVSS.n1671 DVSS.n1670 585
R5986 DVSS.n537 DVSS.n536 585
R5987 DVSS.n1669 DVSS.n537 585
R5988 DVSS.n1667 DVSS.n1666 585
R5989 DVSS.n1668 DVSS.n1667 585
R5990 DVSS.n539 DVSS.n538 585
R5991 DVSS.n1654 DVSS.n538 585
R5992 DVSS.n1657 DVSS.n1656 585
R5993 DVSS.n1656 DVSS.n1655 585
R5994 DVSS.n542 DVSS.n541 585
R5995 DVSS.n543 DVSS.n542 585
R5996 DVSS.n703 DVSS.n702 585
R5997 DVSS.n702 DVSS.n701 585
R5998 DVSS.n711 DVSS.n658 585
R5999 DVSS.n700 DVSS.n658 585
R6000 DVSS.n712 DVSS.n657 585
R6001 DVSS.n699 DVSS.n657 585
R6002 DVSS.n697 DVSS.n656 585
R6003 DVSS.n698 DVSS.n697 585
R6004 DVSS.n719 DVSS.n655 585
R6005 DVSS.n695 DVSS.n655 585
R6006 DVSS.n720 DVSS.n654 585
R6007 DVSS.n694 DVSS.n654 585
R6008 DVSS.n692 DVSS.n653 585
R6009 DVSS.n693 DVSS.n692 585
R6010 DVSS.n724 DVSS.n652 585
R6011 DVSS.n691 DVSS.n652 585
R6012 DVSS.n725 DVSS.n651 585
R6013 DVSS.n690 DVSS.n651 585
R6014 DVSS.n688 DVSS.n650 585
R6015 DVSS.n689 DVSS.n688 585
R6016 DVSS.n729 DVSS.n649 585
R6017 DVSS.n687 DVSS.n649 585
R6018 DVSS.n730 DVSS.n648 585
R6019 DVSS.n686 DVSS.n648 585
R6020 DVSS.n733 DVSS.n647 585
R6021 DVSS.n685 DVSS.n647 585
R6022 DVSS.n734 DVSS.n646 585
R6023 DVSS.n684 DVSS.n646 585
R6024 DVSS.n682 DVSS.n644 585
R6025 DVSS.n683 DVSS.n682 585
R6026 DVSS.n742 DVSS.n643 585
R6027 DVSS.n681 DVSS.n643 585
R6028 DVSS.n743 DVSS.n642 585
R6029 DVSS.n680 DVSS.n642 585
R6030 DVSS.n678 DVSS.n641 585
R6031 DVSS.n679 DVSS.n678 585
R6032 DVSS.n747 DVSS.n640 585
R6033 DVSS.n677 DVSS.n640 585
R6034 DVSS.n748 DVSS.n639 585
R6035 DVSS.n676 DVSS.n639 585
R6036 DVSS.n674 DVSS.n638 585
R6037 DVSS.n675 DVSS.n674 585
R6038 DVSS.n752 DVSS.n637 585
R6039 DVSS.n673 DVSS.n637 585
R6040 DVSS.n753 DVSS.n636 585
R6041 DVSS.n672 DVSS.n636 585
R6042 DVSS.n669 DVSS.n635 585
R6043 DVSS.n670 DVSS.n669 585
R6044 DVSS.n668 DVSS.n662 585
R6045 DVSS.n668 DVSS.n667 585
R6046 DVSS.n659 DVSS.n631 585
R6047 DVSS.n666 DVSS.n659 585
R6048 DVSS.n1332 DVSS.n630 585
R6049 DVSS.n665 DVSS.n630 585
R6050 DVSS.n1333 DVSS.n629 585
R6051 DVSS.n664 DVSS.n629 585
R6052 DVSS.n628 DVSS.n626 585
R6053 DVSS.n663 DVSS.n626 585
R6054 DVSS.n1338 DVSS.n1337 585
R6055 DVSS.n1339 DVSS.n1338 585
R6056 DVSS.n627 DVSS.n625 585
R6057 DVSS.n625 DVSS.n624 585
R6058 DVSS.n1321 DVSS.n1320 585
R6059 DVSS.n1320 DVSS.n1319 585
R6060 DVSS.n759 DVSS.n758 585
R6061 DVSS.n1318 DVSS.n759 585
R6062 DVSS.n1316 DVSS.n1315 585
R6063 DVSS.n1317 DVSS.n1316 585
R6064 DVSS.n762 DVSS.n761 585
R6065 DVSS.n761 DVSS.n760 585
R6066 DVSS.n1310 DVSS.n1309 585
R6067 DVSS.n1309 DVSS.n1308 585
R6068 DVSS.n764 DVSS.n763 585
R6069 DVSS.n1307 DVSS.n764 585
R6070 DVSS.n1305 DVSS.n1304 585
R6071 DVSS.n1306 DVSS.n1305 585
R6072 DVSS.n1300 DVSS.n766 585
R6073 DVSS.n766 DVSS.n765 585
R6074 DVSS.n1299 DVSS.n768 585
R6075 DVSS.n1288 DVSS.n768 585
R6076 DVSS.n773 DVSS.n767 585
R6077 DVSS.n1289 DVSS.n773 585
R6078 DVSS.n1292 DVSS.n1291 585
R6079 DVSS.n1291 DVSS.n1290 585
R6080 DVSS.n772 DVSS.n771 585
R6081 DVSS.n1287 DVSS.n772 585
R6082 DVSS.n1285 DVSS.n1284 585
R6083 DVSS.n1286 DVSS.n1285 585
R6084 DVSS.n776 DVSS.n775 585
R6085 DVSS.n775 DVSS.n774 585
R6086 DVSS.n1279 DVSS.n1278 585
R6087 DVSS.n1278 DVSS.n1277 585
R6088 DVSS.n778 DVSS.n777 585
R6089 DVSS.n1276 DVSS.n778 585
R6090 DVSS.n1274 DVSS.n1273 585
R6091 DVSS.n1275 DVSS.n1274 585
R6092 DVSS.n781 DVSS.n780 585
R6093 DVSS.n780 DVSS.n779 585
R6094 DVSS.n1264 DVSS.n1263 585
R6095 DVSS.n1263 DVSS.n1262 585
R6096 DVSS.n784 DVSS.n783 585
R6097 DVSS.n1150 DVSS.n784 585
R6098 DVSS.n1153 DVSS.n1152 585
R6099 DVSS.n1152 DVSS.n1151 585
R6100 DVSS.n1161 DVSS.n1146 585
R6101 DVSS.n1149 DVSS.n1146 585
R6102 DVSS.n1162 DVSS.n1145 585
R6103 DVSS.n1148 DVSS.n1145 585
R6104 DVSS.n829 DVSS.n827 585
R6105 DVSS.n1147 DVSS.n827 585
R6106 DVSS.n1167 DVSS.n1166 585
R6107 DVSS.n1168 DVSS.n1167 585
R6108 DVSS.n828 DVSS.n826 585
R6109 DVSS.n826 DVSS.n825 585
R6110 DVSS.n1139 DVSS.n1138 585
R6111 DVSS.n1138 DVSS.n1137 585
R6112 DVSS.n831 DVSS.n830 585
R6113 DVSS.n1136 DVSS.n831 585
R6114 DVSS.n1134 DVSS.n1133 585
R6115 DVSS.n1135 DVSS.n1134 585
R6116 DVSS.n834 DVSS.n833 585
R6117 DVSS.n833 DVSS.n832 585
R6118 DVSS.n1128 DVSS.n1127 585
R6119 DVSS.n1127 DVSS.n1126 585
R6120 DVSS.n836 DVSS.n835 585
R6121 DVSS.n1125 DVSS.n836 585
R6122 DVSS.n1123 DVSS.n1122 585
R6123 DVSS.n1124 DVSS.n1123 585
R6124 DVSS.n1118 DVSS.n838 585
R6125 DVSS.n838 DVSS.n837 585
R6126 DVSS.n1117 DVSS.n840 585
R6127 DVSS.n1106 DVSS.n840 585
R6128 DVSS.n845 DVSS.n839 585
R6129 DVSS.n1107 DVSS.n845 585
R6130 DVSS.n1110 DVSS.n1109 585
R6131 DVSS.n1109 DVSS.n1108 585
R6132 DVSS.n844 DVSS.n843 585
R6133 DVSS.n1105 DVSS.n844 585
R6134 DVSS.n1103 DVSS.n1102 585
R6135 DVSS.n1104 DVSS.n1103 585
R6136 DVSS.n848 DVSS.n847 585
R6137 DVSS.n847 DVSS.n846 585
R6138 DVSS.n1097 DVSS.n1096 585
R6139 DVSS.n1096 DVSS.n1095 585
R6140 DVSS.n850 DVSS.n849 585
R6141 DVSS.n1094 DVSS.n850 585
R6142 DVSS.n1092 DVSS.n1091 585
R6143 DVSS.n1093 DVSS.n1092 585
R6144 DVSS.n853 DVSS.n852 585
R6145 DVSS.n852 DVSS.n851 585
R6146 DVSS.n1082 DVSS.n1081 585
R6147 DVSS.n1081 DVSS.n1080 585
R6148 DVSS.n856 DVSS.n855 585
R6149 DVSS.n968 DVSS.n856 585
R6150 DVSS.n971 DVSS.n970 585
R6151 DVSS.n970 DVSS.n969 585
R6152 DVSS.n979 DVSS.n964 585
R6153 DVSS.n967 DVSS.n964 585
R6154 DVSS.n980 DVSS.n963 585
R6155 DVSS.n966 DVSS.n963 585
R6156 DVSS.n901 DVSS.n899 585
R6157 DVSS.n965 DVSS.n899 585
R6158 DVSS.n985 DVSS.n984 585
R6159 DVSS.n986 DVSS.n985 585
R6160 DVSS.n900 DVSS.n898 585
R6161 DVSS.n898 DVSS.n897 585
R6162 DVSS.n957 DVSS.n956 585
R6163 DVSS.n956 DVSS.n955 585
R6164 DVSS.n903 DVSS.n902 585
R6165 DVSS.n923 DVSS.n918 585
R6166 DVSS.n925 DVSS.n924 585
R6167 DVSS.n927 DVSS.n915 585
R6168 DVSS.n929 DVSS.n928 585
R6169 DVSS.n1 DVSS.n0 585
R6170 DVSS.n2605 DVSS.n2602 585
R6171 DVSS.n2606 DVSS.n2600 585
R6172 DVSS.n2599 DVSS.n2596 585
R6173 DVSS.n2597 DVSS.n2590 585
R6174 DVSS.n2613 DVSS.n2589 585
R6175 DVSS.n2614 DVSS.n2587 585
R6176 DVSS.n2586 DVSS.n2583 585
R6177 DVSS.n2584 DVSS.n2576 585
R6178 DVSS.n2622 DVSS.n2575 585
R6179 DVSS.n2623 DVSS.n2573 585
R6180 DVSS.n2572 DVSS.n2570 585
R6181 DVSS.n2572 DVSS.n3 585
R6182 DVSS.n2627 DVSS.n2569 585
R6183 DVSS.n2569 DVSS.n2568 585
R6184 DVSS.n2628 DVSS.n2562 585
R6185 DVSS.n2567 DVSS.n2562 585
R6186 DVSS.n2565 DVSS.n2559 585
R6187 DVSS.n2566 DVSS.n2565 585
R6188 DVSS.n2636 DVSS.n2558 585
R6189 DVSS.n2564 DVSS.n2558 585
R6190 DVSS.n2637 DVSS.n2557 585
R6191 DVSS.n2563 DVSS.n2557 585
R6192 DVSS.n59 DVSS.n57 585
R6193 DVSS.n57 DVSS.n55 585
R6194 DVSS.n2642 DVSS.n2641 585
R6195 DVSS.n2643 DVSS.n2642 585
R6196 DVSS.n58 DVSS.n56 585
R6197 DVSS.n2554 DVSS.n2553 585
R6198 DVSS.n2551 DVSS.n60 585
R6199 DVSS.n2549 DVSS.n2548 585
R6200 DVSS.n62 DVSS.n61 585
R6201 DVSS.n2537 DVSS.n2536 585
R6202 DVSS.n2534 DVSS.n66 585
R6203 DVSS.n2532 DVSS.n2531 585
R6204 DVSS.n68 DVSS.n67 585
R6205 DVSS.n2526 DVSS.n2525 585
R6206 DVSS.n2523 DVSS.n69 585
R6207 DVSS.n2521 DVSS.n2520 585
R6208 DVSS.n71 DVSS.n70 585
R6209 DVSS.n2509 DVSS.n2508 585
R6210 DVSS.n2506 DVSS.n75 585
R6211 DVSS.n2504 DVSS.n2503 585
R6212 DVSS.n77 DVSS.n76 585
R6213 DVSS.n2492 DVSS.n2491 585
R6214 DVSS.n2489 DVSS.n79 585
R6215 DVSS.n2489 DVSS.n53 585
R6216 DVSS.n2488 DVSS.n2487 585
R6217 DVSS.n2488 DVSS.n52 585
R6218 DVSS.n81 DVSS.n80 585
R6219 DVSS.n2474 DVSS.n80 585
R6220 DVSS.n2477 DVSS.n2476 585
R6221 DVSS.n2476 DVSS.n2475 585
R6222 DVSS.n85 DVSS.n84 585
R6223 DVSS.n2473 DVSS.n85 585
R6224 DVSS.n2471 DVSS.n2470 585
R6225 DVSS.n2472 DVSS.n2471 585
R6226 DVSS.n88 DVSS.n87 585
R6227 DVSS.n2462 DVSS.n87 585
R6228 DVSS.n2465 DVSS.n2464 585
R6229 DVSS.n2464 DVSS.n2463 585
R6230 DVSS.n90 DVSS.n89 585
R6231 DVSS.n2458 DVSS.n2457 585
R6232 DVSS.n97 DVSS.n96 585
R6233 DVSS.n2446 DVSS.n2445 585
R6234 DVSS.n2447 DVSS.n2444 585
R6235 DVSS.n2443 DVSS.n105 585
R6236 DVSS.n104 DVSS.n103 585
R6237 DVSS.n2439 DVSS.n2438 585
R6238 DVSS.n2437 DVSS.n106 585
R6239 DVSS.n2435 DVSS.n2434 585
R6240 DVSS.n108 DVSS.n107 585
R6241 DVSS.n2424 DVSS.n2422 585
R6242 DVSS.n2425 DVSS.n2420 585
R6243 DVSS.n2418 DVSS.n114 585
R6244 DVSS.n2417 DVSS.n2416 585
R6245 DVSS.n2405 DVSS.n116 585
R6246 DVSS.n2407 DVSS.n2406 585
R6247 DVSS.n2403 DVSS.n119 585
R6248 DVSS.n2402 DVSS.n2401 585
R6249 DVSS.n2402 DVSS.n92 585
R6250 DVSS.n121 DVSS.n120 585
R6251 DVSS.n2387 DVSS.n120 585
R6252 DVSS.n2390 DVSS.n2389 585
R6253 DVSS.n2389 DVSS.n2388 585
R6254 DVSS.n125 DVSS.n124 585
R6255 DVSS.n2386 DVSS.n125 585
R6256 DVSS.n2384 DVSS.n2383 585
R6257 DVSS.n2385 DVSS.n2384 585
R6258 DVSS.n128 DVSS.n127 585
R6259 DVSS.n127 DVSS.n126 585
R6260 DVSS.n2378 DVSS.n2377 585
R6261 DVSS.n2377 DVSS.n2376 585
R6262 DVSS.n130 DVSS.n129 585
R6263 DVSS.n131 DVSS.n130 585
R6264 DVSS.n2290 DVSS.n2289 585
R6265 DVSS.n299 DVSS.n298 585
R6266 DVSS.n2284 DVSS.n2283 585
R6267 DVSS.n2282 DVSS.n303 585
R6268 DVSS.n302 DVSS.n301 585
R6269 DVSS.n2271 DVSS.n2270 585
R6270 DVSS.n2269 DVSS.n2268 585
R6271 DVSS.n2262 DVSS.n305 585
R6272 DVSS.n2264 DVSS.n2263 585
R6273 DVSS.n2260 DVSS.n306 585
R6274 DVSS.n2259 DVSS.n2258 585
R6275 DVSS.n2248 DVSS.n308 585
R6276 DVSS.n2250 DVSS.n2249 585
R6277 DVSS.n2246 DVSS.n315 585
R6278 DVSS.n2245 DVSS.n2244 585
R6279 DVSS.n2233 DVSS.n317 585
R6280 DVSS.n2235 DVSS.n2234 585
R6281 DVSS.n2231 DVSS.n320 585
R6282 DVSS.n2230 DVSS.n2229 585
R6283 DVSS.n2230 DVSS.n294 585
R6284 DVSS.n322 DVSS.n321 585
R6285 DVSS.n321 DVSS.n293 585
R6286 DVSS.n2218 DVSS.n2217 585
R6287 DVSS.n2217 DVSS.n2216 585
R6288 DVSS.n326 DVSS.n325 585
R6289 DVSS.n2215 DVSS.n326 585
R6290 DVSS.n2213 DVSS.n2212 585
R6291 DVSS.n2214 DVSS.n2213 585
R6292 DVSS.n329 DVSS.n328 585
R6293 DVSS.n328 DVSS.n327 585
R6294 DVSS.n2207 DVSS.n2206 585
R6295 DVSS.n2206 DVSS.n2205 585
R6296 DVSS.n331 DVSS.n330 585
R6297 DVSS.n332 DVSS.n331 585
R6298 DVSS.n2108 DVSS.n2107 585
R6299 DVSS.n371 DVSS.n370 585
R6300 DVSS.n2102 DVSS.n2101 585
R6301 DVSS.n2100 DVSS.n375 585
R6302 DVSS.n374 DVSS.n373 585
R6303 DVSS.n2089 DVSS.n2088 585
R6304 DVSS.n2087 DVSS.n2086 585
R6305 DVSS.n2080 DVSS.n377 585
R6306 DVSS.n2082 DVSS.n2081 585
R6307 DVSS.n2078 DVSS.n378 585
R6308 DVSS.n2077 DVSS.n2076 585
R6309 DVSS.n2066 DVSS.n380 585
R6310 DVSS.n2068 DVSS.n2067 585
R6311 DVSS.n2064 DVSS.n387 585
R6312 DVSS.n2063 DVSS.n2062 585
R6313 DVSS.n2051 DVSS.n389 585
R6314 DVSS.n2053 DVSS.n2052 585
R6315 DVSS.n2049 DVSS.n392 585
R6316 DVSS.n2048 DVSS.n2047 585
R6317 DVSS.n2048 DVSS.n366 585
R6318 DVSS.n394 DVSS.n393 585
R6319 DVSS.n393 DVSS.n365 585
R6320 DVSS.n2036 DVSS.n2035 585
R6321 DVSS.n2035 DVSS.n2034 585
R6322 DVSS.n398 DVSS.n397 585
R6323 DVSS.n2033 DVSS.n398 585
R6324 DVSS.n2031 DVSS.n2030 585
R6325 DVSS.n2032 DVSS.n2031 585
R6326 DVSS.n401 DVSS.n400 585
R6327 DVSS.n400 DVSS.n399 585
R6328 DVSS.n2025 DVSS.n2024 585
R6329 DVSS.n2024 DVSS.n2023 585
R6330 DVSS.n403 DVSS.n402 585
R6331 DVSS.n404 DVSS.n403 585
R6332 DVSS.n1926 DVSS.n1925 585
R6333 DVSS.n443 DVSS.n442 585
R6334 DVSS.n1920 DVSS.n1919 585
R6335 DVSS.n1918 DVSS.n447 585
R6336 DVSS.n446 DVSS.n445 585
R6337 DVSS.n1907 DVSS.n1906 585
R6338 DVSS.n1905 DVSS.n1904 585
R6339 DVSS.n1898 DVSS.n449 585
R6340 DVSS.n1900 DVSS.n1899 585
R6341 DVSS.n1896 DVSS.n450 585
R6342 DVSS.n1895 DVSS.n1894 585
R6343 DVSS.n1884 DVSS.n452 585
R6344 DVSS.n1886 DVSS.n1885 585
R6345 DVSS.n1882 DVSS.n459 585
R6346 DVSS.n1881 DVSS.n1880 585
R6347 DVSS.n1869 DVSS.n461 585
R6348 DVSS.n1871 DVSS.n1870 585
R6349 DVSS.n1867 DVSS.n464 585
R6350 DVSS.n1866 DVSS.n1865 585
R6351 DVSS.n1866 DVSS.n438 585
R6352 DVSS.n466 DVSS.n465 585
R6353 DVSS.n465 DVSS.n437 585
R6354 DVSS.n1854 DVSS.n1853 585
R6355 DVSS.n1853 DVSS.n1852 585
R6356 DVSS.n470 DVSS.n469 585
R6357 DVSS.n1851 DVSS.n470 585
R6358 DVSS.n1849 DVSS.n1848 585
R6359 DVSS.n1850 DVSS.n1849 585
R6360 DVSS.n473 DVSS.n472 585
R6361 DVSS.n472 DVSS.n471 585
R6362 DVSS.n1843 DVSS.n1842 585
R6363 DVSS.n1842 DVSS.n1841 585
R6364 DVSS.n475 DVSS.n474 585
R6365 DVSS.n476 DVSS.n475 585
R6366 DVSS.n1593 DVSS.n1592 585
R6367 DVSS.n1565 DVSS.n1563 585
R6368 DVSS.n1597 DVSS.n1562 585
R6369 DVSS.n1598 DVSS.n1561 585
R6370 DVSS.n1587 DVSS.n1556 585
R6371 DVSS.n1607 DVSS.n1555 585
R6372 DVSS.n1608 DVSS.n1554 585
R6373 DVSS.n1585 DVSS.n1553 585
R6374 DVSS.n1612 DVSS.n1552 585
R6375 DVSS.n1613 DVSS.n1551 585
R6376 DVSS.n1575 DVSS.n1550 585
R6377 DVSS.n1574 DVSS.n1544 585
R6378 DVSS.n1620 DVSS.n1543 585
R6379 DVSS.n1621 DVSS.n1542 585
R6380 DVSS.n1579 DVSS.n1541 585
R6381 DVSS.n1578 DVSS.n1534 585
R6382 DVSS.n1629 DVSS.n1533 585
R6383 DVSS.n1630 DVSS.n1532 585
R6384 DVSS.n1582 DVSS.n1530 585
R6385 DVSS.n1583 DVSS.n1582 585
R6386 DVSS.n1634 DVSS.n1529 585
R6387 DVSS.n1571 DVSS.n1529 585
R6388 DVSS.n1635 DVSS.n1528 585
R6389 DVSS.n1570 DVSS.n1528 585
R6390 DVSS.n1568 DVSS.n1525 585
R6391 DVSS.n1569 DVSS.n1568 585
R6392 DVSS.n1643 DVSS.n1524 585
R6393 DVSS.n1567 DVSS.n1524 585
R6394 DVSS.n1644 DVSS.n1523 585
R6395 DVSS.n1566 DVSS.n1523 585
R6396 DVSS.n551 DVSS.n549 585
R6397 DVSS.n549 DVSS.n547 585
R6398 DVSS.n1649 DVSS.n1648 585
R6399 DVSS.n1650 DVSS.n1649 585
R6400 DVSS.n550 DVSS.n548 585
R6401 DVSS.n1520 DVSS.n1519 585
R6402 DVSS.n1517 DVSS.n552 585
R6403 DVSS.n1515 DVSS.n1514 585
R6404 DVSS.n554 DVSS.n553 585
R6405 DVSS.n1503 DVSS.n1502 585
R6406 DVSS.n1500 DVSS.n558 585
R6407 DVSS.n1498 DVSS.n1497 585
R6408 DVSS.n560 DVSS.n559 585
R6409 DVSS.n1492 DVSS.n1491 585
R6410 DVSS.n1489 DVSS.n561 585
R6411 DVSS.n1487 DVSS.n1486 585
R6412 DVSS.n563 DVSS.n562 585
R6413 DVSS.n1475 DVSS.n1474 585
R6414 DVSS.n1472 DVSS.n567 585
R6415 DVSS.n1470 DVSS.n1469 585
R6416 DVSS.n569 DVSS.n568 585
R6417 DVSS.n1458 DVSS.n1457 585
R6418 DVSS.n1455 DVSS.n571 585
R6419 DVSS.n1455 DVSS.n545 585
R6420 DVSS.n1454 DVSS.n1453 585
R6421 DVSS.n1454 DVSS.n544 585
R6422 DVSS.n573 DVSS.n572 585
R6423 DVSS.n1440 DVSS.n572 585
R6424 DVSS.n1443 DVSS.n1442 585
R6425 DVSS.n1442 DVSS.n1441 585
R6426 DVSS.n577 DVSS.n576 585
R6427 DVSS.n1439 DVSS.n577 585
R6428 DVSS.n1437 DVSS.n1436 585
R6429 DVSS.n1438 DVSS.n1437 585
R6430 DVSS.n580 DVSS.n579 585
R6431 DVSS.n1428 DVSS.n579 585
R6432 DVSS.n1431 DVSS.n1430 585
R6433 DVSS.n1430 DVSS.n1429 585
R6434 DVSS.n582 DVSS.n581 585
R6435 DVSS.n1424 DVSS.n1423 585
R6436 DVSS.n589 DVSS.n588 585
R6437 DVSS.n1412 DVSS.n1411 585
R6438 DVSS.n1413 DVSS.n1410 585
R6439 DVSS.n1409 DVSS.n597 585
R6440 DVSS.n596 DVSS.n595 585
R6441 DVSS.n1405 DVSS.n1404 585
R6442 DVSS.n1403 DVSS.n598 585
R6443 DVSS.n1401 DVSS.n1400 585
R6444 DVSS.n600 DVSS.n599 585
R6445 DVSS.n1390 DVSS.n1388 585
R6446 DVSS.n1391 DVSS.n1386 585
R6447 DVSS.n1384 DVSS.n606 585
R6448 DVSS.n1383 DVSS.n1382 585
R6449 DVSS.n1371 DVSS.n608 585
R6450 DVSS.n1373 DVSS.n1372 585
R6451 DVSS.n1369 DVSS.n611 585
R6452 DVSS.n1368 DVSS.n1367 585
R6453 DVSS.n1368 DVSS.n584 585
R6454 DVSS.n613 DVSS.n612 585
R6455 DVSS.n1353 DVSS.n612 585
R6456 DVSS.n1356 DVSS.n1355 585
R6457 DVSS.n1355 DVSS.n1354 585
R6458 DVSS.n617 DVSS.n616 585
R6459 DVSS.n1352 DVSS.n617 585
R6460 DVSS.n1350 DVSS.n1349 585
R6461 DVSS.n1351 DVSS.n1350 585
R6462 DVSS.n620 DVSS.n619 585
R6463 DVSS.n619 DVSS.n618 585
R6464 DVSS.n1344 DVSS.n1343 585
R6465 DVSS.n1343 DVSS.n1342 585
R6466 DVSS.n622 DVSS.n621 585
R6467 DVSS.n623 DVSS.n622 585
R6468 DVSS.n1256 DVSS.n1255 585
R6469 DVSS.n791 DVSS.n790 585
R6470 DVSS.n1250 DVSS.n1249 585
R6471 DVSS.n1248 DVSS.n795 585
R6472 DVSS.n794 DVSS.n793 585
R6473 DVSS.n1237 DVSS.n1236 585
R6474 DVSS.n1235 DVSS.n1234 585
R6475 DVSS.n1228 DVSS.n797 585
R6476 DVSS.n1230 DVSS.n1229 585
R6477 DVSS.n1226 DVSS.n798 585
R6478 DVSS.n1225 DVSS.n1224 585
R6479 DVSS.n1214 DVSS.n800 585
R6480 DVSS.n1216 DVSS.n1215 585
R6481 DVSS.n1212 DVSS.n807 585
R6482 DVSS.n1211 DVSS.n1210 585
R6483 DVSS.n1199 DVSS.n809 585
R6484 DVSS.n1201 DVSS.n1200 585
R6485 DVSS.n1197 DVSS.n812 585
R6486 DVSS.n1196 DVSS.n1195 585
R6487 DVSS.n1196 DVSS.n786 585
R6488 DVSS.n814 DVSS.n813 585
R6489 DVSS.n813 DVSS.n785 585
R6490 DVSS.n1184 DVSS.n1183 585
R6491 DVSS.n1183 DVSS.n1182 585
R6492 DVSS.n818 DVSS.n817 585
R6493 DVSS.n1181 DVSS.n818 585
R6494 DVSS.n1179 DVSS.n1178 585
R6495 DVSS.n1180 DVSS.n1179 585
R6496 DVSS.n821 DVSS.n820 585
R6497 DVSS.n820 DVSS.n819 585
R6498 DVSS.n1173 DVSS.n1172 585
R6499 DVSS.n1172 DVSS.n1171 585
R6500 DVSS.n823 DVSS.n822 585
R6501 DVSS.n824 DVSS.n823 585
R6502 DVSS.n1074 DVSS.n1073 585
R6503 DVSS.n863 DVSS.n862 585
R6504 DVSS.n1068 DVSS.n1067 585
R6505 DVSS.n1066 DVSS.n867 585
R6506 DVSS.n866 DVSS.n865 585
R6507 DVSS.n1055 DVSS.n1054 585
R6508 DVSS.n1053 DVSS.n1052 585
R6509 DVSS.n1046 DVSS.n869 585
R6510 DVSS.n1048 DVSS.n1047 585
R6511 DVSS.n1044 DVSS.n870 585
R6512 DVSS.n1043 DVSS.n1042 585
R6513 DVSS.n1032 DVSS.n872 585
R6514 DVSS.n1034 DVSS.n1033 585
R6515 DVSS.n1030 DVSS.n879 585
R6516 DVSS.n1029 DVSS.n1028 585
R6517 DVSS.n1017 DVSS.n881 585
R6518 DVSS.n1019 DVSS.n1018 585
R6519 DVSS.n1015 DVSS.n884 585
R6520 DVSS.n1014 DVSS.n1013 585
R6521 DVSS.n1014 DVSS.n858 585
R6522 DVSS.n886 DVSS.n885 585
R6523 DVSS.n885 DVSS.n857 585
R6524 DVSS.n1002 DVSS.n1001 585
R6525 DVSS.n1001 DVSS.n1000 585
R6526 DVSS.n890 DVSS.n889 585
R6527 DVSS.n999 DVSS.n890 585
R6528 DVSS.n997 DVSS.n996 585
R6529 DVSS.n998 DVSS.n997 585
R6530 DVSS.n893 DVSS.n892 585
R6531 DVSS.n892 DVSS.n891 585
R6532 DVSS.n991 DVSS.n990 585
R6533 DVSS.n990 DVSS.n989 585
R6534 DVSS.n895 DVSS.n894 585
R6535 DVSS.n896 DVSS.n895 585
R6536 DVSS.n951 DVSS.n950 585
R6537 DVSS.n908 DVSS.n907 585
R6538 DVSS.n945 DVSS.n944 585
R6539 DVSS.n943 DVSS.n912 585
R6540 DVSS.n911 DVSS.n910 585
R6541 DVSS.t116 DVSS.n857 552.341
R6542 DVSS.t217 DVSS.n785 552.341
R6543 DVSS.t9 DVSS.n1353 552.341
R6544 DVSS.t42 DVSS.n544 552.341
R6545 DVSS.n1571 DVSS.t59 552.341
R6546 DVSS.t205 DVSS.n437 552.341
R6547 DVSS.t257 DVSS.n365 552.341
R6548 DVSS.t84 DVSS.n293 552.341
R6549 DVSS.t255 DVSS.n2387 552.341
R6550 DVSS.t96 DVSS.n52 552.341
R6551 DVSS.n2568 DVSS.t156 552.341
R6552 DVSS.n928 DVSS.n927 539.294
R6553 DVSS.n925 DVSS.n918 539.294
R6554 DVSS.n956 DVSS.n903 539.294
R6555 DVSS.n956 DVSS.n898 539.294
R6556 DVSS.n985 DVSS.n898 539.294
R6557 DVSS.n985 DVSS.n899 539.294
R6558 DVSS.n963 DVSS.n899 539.294
R6559 DVSS.n964 DVSS.n963 539.294
R6560 DVSS.n970 DVSS.n964 539.294
R6561 DVSS.n970 DVSS.n856 539.294
R6562 DVSS.n1081 DVSS.n856 539.294
R6563 DVSS.n1081 DVSS.n852 539.294
R6564 DVSS.n1092 DVSS.n852 539.294
R6565 DVSS.n1092 DVSS.n850 539.294
R6566 DVSS.n1096 DVSS.n850 539.294
R6567 DVSS.n1096 DVSS.n847 539.294
R6568 DVSS.n1103 DVSS.n847 539.294
R6569 DVSS.n1103 DVSS.n844 539.294
R6570 DVSS.n1109 DVSS.n844 539.294
R6571 DVSS.n1109 DVSS.n845 539.294
R6572 DVSS.n845 DVSS.n840 539.294
R6573 DVSS.n840 DVSS.n838 539.294
R6574 DVSS.n1123 DVSS.n838 539.294
R6575 DVSS.n1123 DVSS.n836 539.294
R6576 DVSS.n1127 DVSS.n836 539.294
R6577 DVSS.n1127 DVSS.n833 539.294
R6578 DVSS.n1134 DVSS.n833 539.294
R6579 DVSS.n1134 DVSS.n831 539.294
R6580 DVSS.n1138 DVSS.n831 539.294
R6581 DVSS.n1138 DVSS.n826 539.294
R6582 DVSS.n1167 DVSS.n826 539.294
R6583 DVSS.n1167 DVSS.n827 539.294
R6584 DVSS.n1145 DVSS.n827 539.294
R6585 DVSS.n1146 DVSS.n1145 539.294
R6586 DVSS.n1152 DVSS.n1146 539.294
R6587 DVSS.n1152 DVSS.n784 539.294
R6588 DVSS.n1263 DVSS.n784 539.294
R6589 DVSS.n1263 DVSS.n780 539.294
R6590 DVSS.n1274 DVSS.n780 539.294
R6591 DVSS.n1274 DVSS.n778 539.294
R6592 DVSS.n1278 DVSS.n778 539.294
R6593 DVSS.n1278 DVSS.n775 539.294
R6594 DVSS.n1285 DVSS.n775 539.294
R6595 DVSS.n1285 DVSS.n772 539.294
R6596 DVSS.n1291 DVSS.n772 539.294
R6597 DVSS.n1291 DVSS.n773 539.294
R6598 DVSS.n773 DVSS.n768 539.294
R6599 DVSS.n768 DVSS.n766 539.294
R6600 DVSS.n1305 DVSS.n766 539.294
R6601 DVSS.n1305 DVSS.n764 539.294
R6602 DVSS.n1309 DVSS.n764 539.294
R6603 DVSS.n1309 DVSS.n761 539.294
R6604 DVSS.n1316 DVSS.n761 539.294
R6605 DVSS.n1316 DVSS.n759 539.294
R6606 DVSS.n1320 DVSS.n759 539.294
R6607 DVSS.n1320 DVSS.n625 539.294
R6608 DVSS.n1338 DVSS.n625 539.294
R6609 DVSS.n1338 DVSS.n626 539.294
R6610 DVSS.n629 DVSS.n626 539.294
R6611 DVSS.n630 DVSS.n629 539.294
R6612 DVSS.n659 DVSS.n630 539.294
R6613 DVSS.n668 DVSS.n659 539.294
R6614 DVSS.n669 DVSS.n668 539.294
R6615 DVSS.n669 DVSS.n636 539.294
R6616 DVSS.n637 DVSS.n636 539.294
R6617 DVSS.n674 DVSS.n637 539.294
R6618 DVSS.n674 DVSS.n639 539.294
R6619 DVSS.n640 DVSS.n639 539.294
R6620 DVSS.n678 DVSS.n640 539.294
R6621 DVSS.n678 DVSS.n642 539.294
R6622 DVSS.n643 DVSS.n642 539.294
R6623 DVSS.n682 DVSS.n643 539.294
R6624 DVSS.n682 DVSS.n646 539.294
R6625 DVSS.n647 DVSS.n646 539.294
R6626 DVSS.n648 DVSS.n647 539.294
R6627 DVSS.n649 DVSS.n648 539.294
R6628 DVSS.n688 DVSS.n649 539.294
R6629 DVSS.n688 DVSS.n651 539.294
R6630 DVSS.n652 DVSS.n651 539.294
R6631 DVSS.n692 DVSS.n652 539.294
R6632 DVSS.n692 DVSS.n654 539.294
R6633 DVSS.n655 DVSS.n654 539.294
R6634 DVSS.n697 DVSS.n655 539.294
R6635 DVSS.n697 DVSS.n657 539.294
R6636 DVSS.n658 DVSS.n657 539.294
R6637 DVSS.n702 DVSS.n658 539.294
R6638 DVSS.n702 DVSS.n542 539.294
R6639 DVSS.n1656 DVSS.n542 539.294
R6640 DVSS.n1656 DVSS.n538 539.294
R6641 DVSS.n1667 DVSS.n538 539.294
R6642 DVSS.n1667 DVSS.n537 539.294
R6643 DVSS.n1671 DVSS.n537 539.294
R6644 DVSS.n1671 DVSS.n534 539.294
R6645 DVSS.n1678 DVSS.n534 539.294
R6646 DVSS.n1678 DVSS.n532 539.294
R6647 DVSS.n1683 DVSS.n532 539.294
R6648 DVSS.n1683 DVSS.n529 539.294
R6649 DVSS.n1695 DVSS.n529 539.294
R6650 DVSS.n1695 DVSS.n528 539.294
R6651 DVSS.n1699 DVSS.n528 539.294
R6652 DVSS.n1699 DVSS.n525 539.294
R6653 DVSS.n1706 DVSS.n525 539.294
R6654 DVSS.n1706 DVSS.n523 539.294
R6655 DVSS.n1711 DVSS.n523 539.294
R6656 DVSS.n1711 DVSS.n520 539.294
R6657 DVSS.n1718 DVSS.n520 539.294
R6658 DVSS.n1719 DVSS.n1718 539.294
R6659 DVSS.n1719 DVSS.n514 539.294
R6660 DVSS.n515 DVSS.n514 539.294
R6661 DVSS.n1724 DVSS.n515 539.294
R6662 DVSS.n1724 DVSS.n517 539.294
R6663 DVSS.n1728 DVSS.n517 539.294
R6664 DVSS.n1728 DVSS.n508 539.294
R6665 DVSS.n1751 DVSS.n508 539.294
R6666 DVSS.n1751 DVSS.n506 539.294
R6667 DVSS.n1756 DVSS.n506 539.294
R6668 DVSS.n1756 DVSS.n503 539.294
R6669 DVSS.n1763 DVSS.n503 539.294
R6670 DVSS.n1763 DVSS.n501 539.294
R6671 DVSS.n1767 DVSS.n501 539.294
R6672 DVSS.n1767 DVSS.n498 539.294
R6673 DVSS.n1774 DVSS.n498 539.294
R6674 DVSS.n1774 DVSS.n496 539.294
R6675 DVSS.n1780 DVSS.n496 539.294
R6676 DVSS.n1780 DVSS.n492 539.294
R6677 DVSS.n492 DVSS.n490 539.294
R6678 DVSS.n1793 DVSS.n490 539.294
R6679 DVSS.n1793 DVSS.n488 539.294
R6680 DVSS.n1797 DVSS.n488 539.294
R6681 DVSS.n1797 DVSS.n485 539.294
R6682 DVSS.n1804 DVSS.n485 539.294
R6683 DVSS.n1804 DVSS.n483 539.294
R6684 DVSS.n1808 DVSS.n483 539.294
R6685 DVSS.n1808 DVSS.n478 539.294
R6686 DVSS.n1837 DVSS.n478 539.294
R6687 DVSS.n1837 DVSS.n479 539.294
R6688 DVSS.n1815 DVSS.n479 539.294
R6689 DVSS.n1816 DVSS.n1815 539.294
R6690 DVSS.n1822 DVSS.n1816 539.294
R6691 DVSS.n1822 DVSS.n436 539.294
R6692 DVSS.n1933 DVSS.n436 539.294
R6693 DVSS.n1933 DVSS.n432 539.294
R6694 DVSS.n1944 DVSS.n432 539.294
R6695 DVSS.n1944 DVSS.n430 539.294
R6696 DVSS.n1948 DVSS.n430 539.294
R6697 DVSS.n1948 DVSS.n427 539.294
R6698 DVSS.n1955 DVSS.n427 539.294
R6699 DVSS.n1955 DVSS.n424 539.294
R6700 DVSS.n1961 DVSS.n424 539.294
R6701 DVSS.n1961 DVSS.n425 539.294
R6702 DVSS.n425 DVSS.n420 539.294
R6703 DVSS.n420 DVSS.n418 539.294
R6704 DVSS.n1975 DVSS.n418 539.294
R6705 DVSS.n1975 DVSS.n416 539.294
R6706 DVSS.n1979 DVSS.n416 539.294
R6707 DVSS.n1979 DVSS.n413 539.294
R6708 DVSS.n1986 DVSS.n413 539.294
R6709 DVSS.n1986 DVSS.n411 539.294
R6710 DVSS.n1990 DVSS.n411 539.294
R6711 DVSS.n1990 DVSS.n406 539.294
R6712 DVSS.n2019 DVSS.n406 539.294
R6713 DVSS.n2019 DVSS.n407 539.294
R6714 DVSS.n1997 DVSS.n407 539.294
R6715 DVSS.n1998 DVSS.n1997 539.294
R6716 DVSS.n2004 DVSS.n1998 539.294
R6717 DVSS.n2004 DVSS.n364 539.294
R6718 DVSS.n2115 DVSS.n364 539.294
R6719 DVSS.n2115 DVSS.n360 539.294
R6720 DVSS.n2126 DVSS.n360 539.294
R6721 DVSS.n2126 DVSS.n358 539.294
R6722 DVSS.n2130 DVSS.n358 539.294
R6723 DVSS.n2130 DVSS.n355 539.294
R6724 DVSS.n2137 DVSS.n355 539.294
R6725 DVSS.n2137 DVSS.n352 539.294
R6726 DVSS.n2143 DVSS.n352 539.294
R6727 DVSS.n2143 DVSS.n353 539.294
R6728 DVSS.n353 DVSS.n348 539.294
R6729 DVSS.n348 DVSS.n346 539.294
R6730 DVSS.n2157 DVSS.n346 539.294
R6731 DVSS.n2157 DVSS.n344 539.294
R6732 DVSS.n2161 DVSS.n344 539.294
R6733 DVSS.n2161 DVSS.n341 539.294
R6734 DVSS.n2168 DVSS.n341 539.294
R6735 DVSS.n2168 DVSS.n339 539.294
R6736 DVSS.n2172 DVSS.n339 539.294
R6737 DVSS.n2172 DVSS.n334 539.294
R6738 DVSS.n2201 DVSS.n334 539.294
R6739 DVSS.n2201 DVSS.n335 539.294
R6740 DVSS.n2179 DVSS.n335 539.294
R6741 DVSS.n2180 DVSS.n2179 539.294
R6742 DVSS.n2186 DVSS.n2180 539.294
R6743 DVSS.n2186 DVSS.n292 539.294
R6744 DVSS.n2297 DVSS.n292 539.294
R6745 DVSS.n2297 DVSS.n288 539.294
R6746 DVSS.n2308 DVSS.n288 539.294
R6747 DVSS.n2308 DVSS.n286 539.294
R6748 DVSS.n2312 DVSS.n286 539.294
R6749 DVSS.n2312 DVSS.n283 539.294
R6750 DVSS.n2319 DVSS.n283 539.294
R6751 DVSS.n2319 DVSS.n280 539.294
R6752 DVSS.n2325 DVSS.n280 539.294
R6753 DVSS.n2325 DVSS.n281 539.294
R6754 DVSS.n281 DVSS.n276 539.294
R6755 DVSS.n276 DVSS.n274 539.294
R6756 DVSS.n2339 DVSS.n274 539.294
R6757 DVSS.n2339 DVSS.n272 539.294
R6758 DVSS.n2343 DVSS.n272 539.294
R6759 DVSS.n2343 DVSS.n269 539.294
R6760 DVSS.n2350 DVSS.n269 539.294
R6761 DVSS.n2350 DVSS.n267 539.294
R6762 DVSS.n2354 DVSS.n267 539.294
R6763 DVSS.n2354 DVSS.n133 539.294
R6764 DVSS.n2372 DVSS.n133 539.294
R6765 DVSS.n2372 DVSS.n134 539.294
R6766 DVSS.n137 DVSS.n134 539.294
R6767 DVSS.n138 DVSS.n137 539.294
R6768 DVSS.n167 DVSS.n138 539.294
R6769 DVSS.n176 DVSS.n167 539.294
R6770 DVSS.n177 DVSS.n176 539.294
R6771 DVSS.n177 DVSS.n144 539.294
R6772 DVSS.n145 DVSS.n144 539.294
R6773 DVSS.n182 DVSS.n145 539.294
R6774 DVSS.n182 DVSS.n147 539.294
R6775 DVSS.n148 DVSS.n147 539.294
R6776 DVSS.n186 DVSS.n148 539.294
R6777 DVSS.n186 DVSS.n150 539.294
R6778 DVSS.n151 DVSS.n150 539.294
R6779 DVSS.n190 DVSS.n151 539.294
R6780 DVSS.n190 DVSS.n154 539.294
R6781 DVSS.n155 DVSS.n154 539.294
R6782 DVSS.n156 DVSS.n155 539.294
R6783 DVSS.n157 DVSS.n156 539.294
R6784 DVSS.n196 DVSS.n157 539.294
R6785 DVSS.n196 DVSS.n159 539.294
R6786 DVSS.n160 DVSS.n159 539.294
R6787 DVSS.n200 DVSS.n160 539.294
R6788 DVSS.n200 DVSS.n162 539.294
R6789 DVSS.n163 DVSS.n162 539.294
R6790 DVSS.n205 DVSS.n163 539.294
R6791 DVSS.n205 DVSS.n165 539.294
R6792 DVSS.n166 DVSS.n165 539.294
R6793 DVSS.n210 DVSS.n166 539.294
R6794 DVSS.n210 DVSS.n50 539.294
R6795 DVSS.n2649 DVSS.n50 539.294
R6796 DVSS.n2649 DVSS.n46 539.294
R6797 DVSS.n2660 DVSS.n46 539.294
R6798 DVSS.n2660 DVSS.n45 539.294
R6799 DVSS.n2664 DVSS.n45 539.294
R6800 DVSS.n2664 DVSS.n42 539.294
R6801 DVSS.n2671 DVSS.n42 539.294
R6802 DVSS.n2671 DVSS.n40 539.294
R6803 DVSS.n2676 DVSS.n40 539.294
R6804 DVSS.n2676 DVSS.n37 539.294
R6805 DVSS.n2688 DVSS.n37 539.294
R6806 DVSS.n2688 DVSS.n36 539.294
R6807 DVSS.n2692 DVSS.n36 539.294
R6808 DVSS.n2692 DVSS.n33 539.294
R6809 DVSS.n2699 DVSS.n33 539.294
R6810 DVSS.n2699 DVSS.n31 539.294
R6811 DVSS.n2704 DVSS.n31 539.294
R6812 DVSS.n2704 DVSS.n28 539.294
R6813 DVSS.n2711 DVSS.n28 539.294
R6814 DVSS.n2712 DVSS.n2711 539.294
R6815 DVSS.n2712 DVSS.n22 539.294
R6816 DVSS.n23 DVSS.n22 539.294
R6817 DVSS.n2717 DVSS.n23 539.294
R6818 DVSS.n2717 DVSS.n25 539.294
R6819 DVSS.n2721 DVSS.n25 539.294
R6820 DVSS.n2721 DVSS.n16 539.294
R6821 DVSS.n2744 DVSS.n16 539.294
R6822 DVSS.n2744 DVSS.n14 539.294
R6823 DVSS.n2749 DVSS.n14 539.294
R6824 DVSS.n2749 DVSS.n9 539.294
R6825 DVSS.n2782 DVSS.n9 539.294
R6826 DVSS.n2782 DVSS.n10 539.294
R6827 DVSS.n2754 DVSS.n2753 539.294
R6828 DVSS.n2757 DVSS.n2756 539.294
R6829 DVSS.n2759 DVSS.n2758 539.294
R6830 DVSS.n912 DVSS.n911 539.294
R6831 DVSS.n944 DVSS.n907 539.294
R6832 DVSS.n951 DVSS.n895 539.294
R6833 DVSS.n990 DVSS.n895 539.294
R6834 DVSS.n990 DVSS.n892 539.294
R6835 DVSS.n997 DVSS.n892 539.294
R6836 DVSS.n997 DVSS.n890 539.294
R6837 DVSS.n1001 DVSS.n890 539.294
R6838 DVSS.n1001 DVSS.n885 539.294
R6839 DVSS.n1014 DVSS.n885 539.294
R6840 DVSS.n1015 DVSS.n1014 539.294
R6841 DVSS.n1018 DVSS.n1017 539.294
R6842 DVSS.n1030 DVSS.n1029 539.294
R6843 DVSS.n1033 DVSS.n1032 539.294
R6844 DVSS.n1044 DVSS.n1043 539.294
R6845 DVSS.n1047 DVSS.n1046 539.294
R6846 DVSS.n1054 DVSS.n1053 539.294
R6847 DVSS.n867 DVSS.n866 539.294
R6848 DVSS.n1067 DVSS.n862 539.294
R6849 DVSS.n1074 DVSS.n823 539.294
R6850 DVSS.n1172 DVSS.n823 539.294
R6851 DVSS.n1172 DVSS.n820 539.294
R6852 DVSS.n1179 DVSS.n820 539.294
R6853 DVSS.n1179 DVSS.n818 539.294
R6854 DVSS.n1183 DVSS.n818 539.294
R6855 DVSS.n1183 DVSS.n813 539.294
R6856 DVSS.n1196 DVSS.n813 539.294
R6857 DVSS.n1197 DVSS.n1196 539.294
R6858 DVSS.n1200 DVSS.n1199 539.294
R6859 DVSS.n1212 DVSS.n1211 539.294
R6860 DVSS.n1215 DVSS.n1214 539.294
R6861 DVSS.n1226 DVSS.n1225 539.294
R6862 DVSS.n1229 DVSS.n1228 539.294
R6863 DVSS.n1236 DVSS.n1235 539.294
R6864 DVSS.n795 DVSS.n794 539.294
R6865 DVSS.n1249 DVSS.n790 539.294
R6866 DVSS.n1256 DVSS.n622 539.294
R6867 DVSS.n1343 DVSS.n622 539.294
R6868 DVSS.n1343 DVSS.n619 539.294
R6869 DVSS.n1350 DVSS.n619 539.294
R6870 DVSS.n1350 DVSS.n617 539.294
R6871 DVSS.n1355 DVSS.n617 539.294
R6872 DVSS.n1355 DVSS.n612 539.294
R6873 DVSS.n1368 DVSS.n612 539.294
R6874 DVSS.n1369 DVSS.n1368 539.294
R6875 DVSS.n1372 DVSS.n1371 539.294
R6876 DVSS.n1384 DVSS.n1383 539.294
R6877 DVSS.n1388 DVSS.n1386 539.294
R6878 DVSS.n1401 DVSS.n599 539.294
R6879 DVSS.n1404 DVSS.n1403 539.294
R6880 DVSS.n597 DVSS.n596 539.294
R6881 DVSS.n1411 DVSS.n1410 539.294
R6882 DVSS.n1424 DVSS.n588 539.294
R6883 DVSS.n1430 DVSS.n582 539.294
R6884 DVSS.n1430 DVSS.n579 539.294
R6885 DVSS.n1437 DVSS.n579 539.294
R6886 DVSS.n1437 DVSS.n577 539.294
R6887 DVSS.n1442 DVSS.n577 539.294
R6888 DVSS.n1442 DVSS.n572 539.294
R6889 DVSS.n1454 DVSS.n572 539.294
R6890 DVSS.n1455 DVSS.n1454 539.294
R6891 DVSS.n1457 DVSS.n1455 539.294
R6892 DVSS.n1470 DVSS.n568 539.294
R6893 DVSS.n1474 DVSS.n1472 539.294
R6894 DVSS.n1487 DVSS.n562 539.294
R6895 DVSS.n1491 DVSS.n1489 539.294
R6896 DVSS.n1498 DVSS.n559 539.294
R6897 DVSS.n1502 DVSS.n1500 539.294
R6898 DVSS.n1515 DVSS.n553 539.294
R6899 DVSS.n1519 DVSS.n1517 539.294
R6900 DVSS.n1649 DVSS.n548 539.294
R6901 DVSS.n1649 DVSS.n549 539.294
R6902 DVSS.n1523 DVSS.n549 539.294
R6903 DVSS.n1524 DVSS.n1523 539.294
R6904 DVSS.n1568 DVSS.n1524 539.294
R6905 DVSS.n1568 DVSS.n1528 539.294
R6906 DVSS.n1529 DVSS.n1528 539.294
R6907 DVSS.n1582 DVSS.n1529 539.294
R6908 DVSS.n1582 DVSS.n1532 539.294
R6909 DVSS.n1578 DVSS.n1533 539.294
R6910 DVSS.n1579 DVSS.n1542 539.294
R6911 DVSS.n1574 DVSS.n1543 539.294
R6912 DVSS.n1575 DVSS.n1551 539.294
R6913 DVSS.n1585 DVSS.n1552 539.294
R6914 DVSS.n1555 DVSS.n1554 539.294
R6915 DVSS.n1587 DVSS.n1561 539.294
R6916 DVSS.n1565 DVSS.n1562 539.294
R6917 DVSS.n1592 DVSS.n475 539.294
R6918 DVSS.n1842 DVSS.n475 539.294
R6919 DVSS.n1842 DVSS.n472 539.294
R6920 DVSS.n1849 DVSS.n472 539.294
R6921 DVSS.n1849 DVSS.n470 539.294
R6922 DVSS.n1853 DVSS.n470 539.294
R6923 DVSS.n1853 DVSS.n465 539.294
R6924 DVSS.n1866 DVSS.n465 539.294
R6925 DVSS.n1867 DVSS.n1866 539.294
R6926 DVSS.n1870 DVSS.n1869 539.294
R6927 DVSS.n1882 DVSS.n1881 539.294
R6928 DVSS.n1885 DVSS.n1884 539.294
R6929 DVSS.n1896 DVSS.n1895 539.294
R6930 DVSS.n1899 DVSS.n1898 539.294
R6931 DVSS.n1906 DVSS.n1905 539.294
R6932 DVSS.n447 DVSS.n446 539.294
R6933 DVSS.n1919 DVSS.n442 539.294
R6934 DVSS.n1926 DVSS.n403 539.294
R6935 DVSS.n2024 DVSS.n403 539.294
R6936 DVSS.n2024 DVSS.n400 539.294
R6937 DVSS.n2031 DVSS.n400 539.294
R6938 DVSS.n2031 DVSS.n398 539.294
R6939 DVSS.n2035 DVSS.n398 539.294
R6940 DVSS.n2035 DVSS.n393 539.294
R6941 DVSS.n2048 DVSS.n393 539.294
R6942 DVSS.n2049 DVSS.n2048 539.294
R6943 DVSS.n2052 DVSS.n2051 539.294
R6944 DVSS.n2064 DVSS.n2063 539.294
R6945 DVSS.n2067 DVSS.n2066 539.294
R6946 DVSS.n2078 DVSS.n2077 539.294
R6947 DVSS.n2081 DVSS.n2080 539.294
R6948 DVSS.n2088 DVSS.n2087 539.294
R6949 DVSS.n375 DVSS.n374 539.294
R6950 DVSS.n2101 DVSS.n370 539.294
R6951 DVSS.n2108 DVSS.n331 539.294
R6952 DVSS.n2206 DVSS.n331 539.294
R6953 DVSS.n2206 DVSS.n328 539.294
R6954 DVSS.n2213 DVSS.n328 539.294
R6955 DVSS.n2213 DVSS.n326 539.294
R6956 DVSS.n2217 DVSS.n326 539.294
R6957 DVSS.n2217 DVSS.n321 539.294
R6958 DVSS.n2230 DVSS.n321 539.294
R6959 DVSS.n2231 DVSS.n2230 539.294
R6960 DVSS.n2234 DVSS.n2233 539.294
R6961 DVSS.n2246 DVSS.n2245 539.294
R6962 DVSS.n2249 DVSS.n2248 539.294
R6963 DVSS.n2260 DVSS.n2259 539.294
R6964 DVSS.n2263 DVSS.n2262 539.294
R6965 DVSS.n2270 DVSS.n2269 539.294
R6966 DVSS.n303 DVSS.n302 539.294
R6967 DVSS.n2283 DVSS.n298 539.294
R6968 DVSS.n2290 DVSS.n130 539.294
R6969 DVSS.n2377 DVSS.n130 539.294
R6970 DVSS.n2377 DVSS.n127 539.294
R6971 DVSS.n2384 DVSS.n127 539.294
R6972 DVSS.n2384 DVSS.n125 539.294
R6973 DVSS.n2389 DVSS.n125 539.294
R6974 DVSS.n2389 DVSS.n120 539.294
R6975 DVSS.n2402 DVSS.n120 539.294
R6976 DVSS.n2403 DVSS.n2402 539.294
R6977 DVSS.n2406 DVSS.n2405 539.294
R6978 DVSS.n2418 DVSS.n2417 539.294
R6979 DVSS.n2422 DVSS.n2420 539.294
R6980 DVSS.n2435 DVSS.n107 539.294
R6981 DVSS.n2438 DVSS.n2437 539.294
R6982 DVSS.n105 DVSS.n104 539.294
R6983 DVSS.n2445 DVSS.n2444 539.294
R6984 DVSS.n2458 DVSS.n96 539.294
R6985 DVSS.n2464 DVSS.n90 539.294
R6986 DVSS.n2464 DVSS.n87 539.294
R6987 DVSS.n2471 DVSS.n87 539.294
R6988 DVSS.n2471 DVSS.n85 539.294
R6989 DVSS.n2476 DVSS.n85 539.294
R6990 DVSS.n2476 DVSS.n80 539.294
R6991 DVSS.n2488 DVSS.n80 539.294
R6992 DVSS.n2489 DVSS.n2488 539.294
R6993 DVSS.n2491 DVSS.n2489 539.294
R6994 DVSS.n2504 DVSS.n76 539.294
R6995 DVSS.n2508 DVSS.n2506 539.294
R6996 DVSS.n2521 DVSS.n70 539.294
R6997 DVSS.n2525 DVSS.n2523 539.294
R6998 DVSS.n2532 DVSS.n67 539.294
R6999 DVSS.n2536 DVSS.n2534 539.294
R7000 DVSS.n2549 DVSS.n61 539.294
R7001 DVSS.n2553 DVSS.n2551 539.294
R7002 DVSS.n2642 DVSS.n56 539.294
R7003 DVSS.n2642 DVSS.n57 539.294
R7004 DVSS.n2557 DVSS.n57 539.294
R7005 DVSS.n2558 DVSS.n2557 539.294
R7006 DVSS.n2565 DVSS.n2558 539.294
R7007 DVSS.n2565 DVSS.n2562 539.294
R7008 DVSS.n2569 DVSS.n2562 539.294
R7009 DVSS.n2572 DVSS.n2569 539.294
R7010 DVSS.n2573 DVSS.n2572 539.294
R7011 DVSS.n2584 DVSS.n2575 539.294
R7012 DVSS.n2587 DVSS.n2586 539.294
R7013 DVSS.n2597 DVSS.n2589 539.294
R7014 DVSS.n2600 DVSS.n2599 539.294
R7015 DVSS.n2602 DVSS.n1 539.294
R7016 DVSS.n1095 DVSS.n1094 526.028
R7017 DVSS.n1095 DVSS.n846 526.028
R7018 DVSS.n1104 DVSS.n846 526.028
R7019 DVSS.n1105 DVSS.n1104 526.028
R7020 DVSS.n1108 DVSS.n1105 526.028
R7021 DVSS.n1107 DVSS.n1106 526.028
R7022 DVSS.n1124 DVSS.n837 526.028
R7023 DVSS.n1125 DVSS.n1124 526.028
R7024 DVSS.n1126 DVSS.n1125 526.028
R7025 DVSS.n1135 DVSS.n832 526.028
R7026 DVSS.n1136 DVSS.n1135 526.028
R7027 DVSS.n1277 DVSS.n1276 526.028
R7028 DVSS.n1277 DVSS.n774 526.028
R7029 DVSS.n1286 DVSS.n774 526.028
R7030 DVSS.n1287 DVSS.n1286 526.028
R7031 DVSS.n1290 DVSS.n1287 526.028
R7032 DVSS.n1289 DVSS.n1288 526.028
R7033 DVSS.n1306 DVSS.n765 526.028
R7034 DVSS.n1307 DVSS.n1306 526.028
R7035 DVSS.n1308 DVSS.n1307 526.028
R7036 DVSS.n1317 DVSS.n760 526.028
R7037 DVSS.n1318 DVSS.n1317 526.028
R7038 DVSS.n676 DVSS.n675 526.028
R7039 DVSS.n677 DVSS.n676 526.028
R7040 DVSS.n679 DVSS.n677 526.028
R7041 DVSS.n680 DVSS.n679 526.028
R7042 DVSS.n681 DVSS.n680 526.028
R7043 DVSS.n684 DVSS.n683 526.028
R7044 DVSS.n686 DVSS.n685 526.028
R7045 DVSS.n687 DVSS.n686 526.028
R7046 DVSS.n689 DVSS.n687 526.028
R7047 DVSS.n691 DVSS.n690 526.028
R7048 DVSS.n693 DVSS.n691 526.028
R7049 DVSS.n1670 DVSS.n533 526.028
R7050 DVSS.n1679 DVSS.n533 526.028
R7051 DVSS.n1680 DVSS.n1679 526.028
R7052 DVSS.n1682 DVSS.n1680 526.028
R7053 DVSS.n1682 DVSS.n1681 526.028
R7054 DVSS.n1697 DVSS.n1696 526.028
R7055 DVSS.n1698 DVSS.n524 526.028
R7056 DVSS.n1707 DVSS.n524 526.028
R7057 DVSS.n1708 DVSS.n1707 526.028
R7058 DVSS.n1710 DVSS.n1709 526.028
R7059 DVSS.n1709 DVSS.n519 526.028
R7060 DVSS.n2663 DVSS.n41 526.028
R7061 DVSS.n2672 DVSS.n41 526.028
R7062 DVSS.n2673 DVSS.n2672 526.028
R7063 DVSS.n2675 DVSS.n2673 526.028
R7064 DVSS.n2675 DVSS.n2674 526.028
R7065 DVSS.n2690 DVSS.n2689 526.028
R7066 DVSS.n2691 DVSS.n32 526.028
R7067 DVSS.n2700 DVSS.n32 526.028
R7068 DVSS.n2701 DVSS.n2700 526.028
R7069 DVSS.n2703 DVSS.n2702 526.028
R7070 DVSS.n2702 DVSS.n27 526.028
R7071 DVSS.n184 DVSS.n183 526.028
R7072 DVSS.n185 DVSS.n184 526.028
R7073 DVSS.n187 DVSS.n185 526.028
R7074 DVSS.n188 DVSS.n187 526.028
R7075 DVSS.n189 DVSS.n188 526.028
R7076 DVSS.n192 DVSS.n191 526.028
R7077 DVSS.n194 DVSS.n193 526.028
R7078 DVSS.n195 DVSS.n194 526.028
R7079 DVSS.n197 DVSS.n195 526.028
R7080 DVSS.n199 DVSS.n198 526.028
R7081 DVSS.n201 DVSS.n199 526.028
R7082 DVSS.n2311 DVSS.n2310 526.028
R7083 DVSS.n2311 DVSS.n282 526.028
R7084 DVSS.n2320 DVSS.n282 526.028
R7085 DVSS.n2321 DVSS.n2320 526.028
R7086 DVSS.n2324 DVSS.n2321 526.028
R7087 DVSS.n2323 DVSS.n2322 526.028
R7088 DVSS.n2340 DVSS.n273 526.028
R7089 DVSS.n2341 DVSS.n2340 526.028
R7090 DVSS.n2342 DVSS.n2341 526.028
R7091 DVSS.n2351 DVSS.n268 526.028
R7092 DVSS.n2352 DVSS.n2351 526.028
R7093 DVSS.n2129 DVSS.n2128 526.028
R7094 DVSS.n2129 DVSS.n354 526.028
R7095 DVSS.n2138 DVSS.n354 526.028
R7096 DVSS.n2139 DVSS.n2138 526.028
R7097 DVSS.n2142 DVSS.n2139 526.028
R7098 DVSS.n2141 DVSS.n2140 526.028
R7099 DVSS.n2158 DVSS.n345 526.028
R7100 DVSS.n2159 DVSS.n2158 526.028
R7101 DVSS.n2160 DVSS.n2159 526.028
R7102 DVSS.n2169 DVSS.n340 526.028
R7103 DVSS.n2170 DVSS.n2169 526.028
R7104 DVSS.n1947 DVSS.n1946 526.028
R7105 DVSS.n1947 DVSS.n426 526.028
R7106 DVSS.n1956 DVSS.n426 526.028
R7107 DVSS.n1957 DVSS.n1956 526.028
R7108 DVSS.n1960 DVSS.n1957 526.028
R7109 DVSS.n1959 DVSS.n1958 526.028
R7110 DVSS.n1976 DVSS.n417 526.028
R7111 DVSS.n1977 DVSS.n1976 526.028
R7112 DVSS.n1978 DVSS.n1977 526.028
R7113 DVSS.n1987 DVSS.n412 526.028
R7114 DVSS.n1988 DVSS.n1987 526.028
R7115 DVSS.n1765 DVSS.n1764 526.028
R7116 DVSS.n1766 DVSS.n1765 526.028
R7117 DVSS.n1766 DVSS.n497 526.028
R7118 DVSS.n1775 DVSS.n497 526.028
R7119 DVSS.n1776 DVSS.n1775 526.028
R7120 DVSS.n1794 DVSS.n489 526.028
R7121 DVSS.n1795 DVSS.n1794 526.028
R7122 DVSS.n1796 DVSS.n1795 526.028
R7123 DVSS.n1805 DVSS.n484 526.028
R7124 DVSS.n1806 DVSS.n1805 526.028
R7125 DVSS.n1078 DVSS.n857 477.447
R7126 DVSS.n1260 DVSS.n785 477.447
R7127 DVSS.n1353 DVSS.n583 477.447
R7128 DVSS.n1652 DVSS.n544 477.447
R7129 DVSS.n1572 DVSS.n1571 477.447
R7130 DVSS.n1930 DVSS.n437 477.447
R7131 DVSS.n2112 DVSS.n365 477.447
R7132 DVSS.n2294 DVSS.n293 477.447
R7133 DVSS.n2387 DVSS.n91 477.447
R7134 DVSS.n2645 DVSS.n52 477.447
R7135 DVSS.n2568 DVSS.n2 477.447
R7136 DVSS.t112 DVSS.n837 465.753
R7137 DVSS.t190 DVSS.n765 465.753
R7138 DVSS.n685 DVSS.t28 465.753
R7139 DVSS.n1698 DVSS.t30 465.753
R7140 DVSS.n2691 DVSS.t72 465.753
R7141 DVSS.n193 DVSS.t227 465.753
R7142 DVSS.t192 DVSS.n273 465.753
R7143 DVSS.t4 DVSS.n345 465.753
R7144 DVSS.t144 DVSS.n417 465.753
R7145 DVSS.t109 DVSS.n489 465.753
R7146 DVSS.n1000 DVSS.t270 458.724
R7147 DVSS.n1182 DVSS.t135 458.724
R7148 DVSS.n1354 DVSS.t0 458.724
R7149 DVSS.t54 DVSS.n1440 458.724
R7150 DVSS.n1570 DVSS.t69 458.724
R7151 DVSS.n1852 DVSS.t48 458.724
R7152 DVSS.n2034 DVSS.t33 458.724
R7153 DVSS.n2216 DVSS.t133 458.724
R7154 DVSS.n2388 DVSS.t50 458.724
R7155 DVSS.t19 DVSS.n2474 458.724
R7156 DVSS.n2567 DVSS.t168 458.724
R7157 DVSS.t270 DVSS.n999 440
R7158 DVSS.t135 DVSS.n1181 440
R7159 DVSS.t0 DVSS.n1352 440
R7160 DVSS.n1441 DVSS.t54 440
R7161 DVSS.t69 DVSS.n1569 440
R7162 DVSS.t48 DVSS.n1851 440
R7163 DVSS.t33 DVSS.n2033 440
R7164 DVSS.t133 DVSS.n2215 440
R7165 DVSS.t50 DVSS.n2386 440
R7166 DVSS.n2475 DVSS.t19 440
R7167 DVSS.t168 DVSS.n2566 440
R7168 DVSS.n1094 DVSS.n1093 406.844
R7169 DVSS.n1276 DVSS.n1275 406.844
R7170 DVSS.n675 DVSS.n673 406.844
R7171 DVSS.n1670 DVSS.n1669 406.844
R7172 DVSS.n1764 DVSS.n502 406.844
R7173 DVSS.n2663 DVSS.n2662 406.844
R7174 DVSS.n183 DVSS.n181 406.844
R7175 DVSS.n2310 DVSS.n2309 406.844
R7176 DVSS.n2128 DVSS.n2127 406.844
R7177 DVSS.n1946 DVSS.n1945 406.844
R7178 DVSS.n1779 DVSS.n1778 394.522
R7179 DVSS.n1137 DVSS.n1136 383.719
R7180 DVSS.n1319 DVSS.n1318 383.719
R7181 DVSS.n694 DVSS.n693 383.719
R7182 DVSS.n1720 DVSS.n519 383.719
R7183 DVSS.n2713 DVSS.n27 383.719
R7184 DVSS.n202 DVSS.n201 383.719
R7185 DVSS.n2353 DVSS.n2352 383.719
R7186 DVSS.n2171 DVSS.n2170 383.719
R7187 DVSS.n1989 DVSS.n1988 383.719
R7188 DVSS.n1807 DVSS.n1806 383.719
R7189 DVSS.t170 DVSS.n1078 358.281
R7190 DVSS.t196 DVSS.n1260 358.281
R7191 DVSS.t146 DVSS.n583 358.281
R7192 DVSS.t229 DVSS.n1652 358.281
R7193 DVSS.n1572 DVSS.t176 358.281
R7194 DVSS.t237 DVSS.n1930 358.281
R7195 DVSS.t182 DVSS.n2112 358.281
R7196 DVSS.t138 DVSS.n2294 358.281
R7197 DVSS.t126 DVSS.n91 358.281
R7198 DVSS.t88 DVSS.n2645 358.281
R7199 DVSS.t22 DVSS.n2 358.281
R7200 DVSS.n955 DVSS.n897 355.257
R7201 DVSS.n967 DVSS.n966 355.257
R7202 DVSS.n969 DVSS.n968 355.257
R7203 DVSS.n1093 DVSS.n851 355.257
R7204 DVSS.n1137 DVSS.n825 355.257
R7205 DVSS.n1149 DVSS.n1148 355.257
R7206 DVSS.n1151 DVSS.n1150 355.257
R7207 DVSS.n1275 DVSS.n779 355.257
R7208 DVSS.n1319 DVSS.n624 355.257
R7209 DVSS.n665 DVSS.n664 355.257
R7210 DVSS.n667 DVSS.n666 355.257
R7211 DVSS.n673 DVSS.n672 355.257
R7212 DVSS.n695 DVSS.n694 355.257
R7213 DVSS.n701 DVSS.n700 355.257
R7214 DVSS.n1655 DVSS.n543 355.257
R7215 DVSS.n1669 DVSS.n1668 355.257
R7216 DVSS.n1721 DVSS.n1720 355.257
R7217 DVSS.n1727 DVSS.n1726 355.257
R7218 DVSS.n1752 DVSS.n507 355.257
R7219 DVSS.n1755 DVSS.n502 355.257
R7220 DVSS.n2714 DVSS.n2713 355.257
R7221 DVSS.n2720 DVSS.n2719 355.257
R7222 DVSS.n2745 DVSS.n15 355.257
R7223 DVSS.n2748 DVSS.n4 355.257
R7224 DVSS.n203 DVSS.n202 355.257
R7225 DVSS.n209 DVSS.n208 355.257
R7226 DVSS.n2648 DVSS.n51 355.257
R7227 DVSS.n2662 DVSS.n2661 355.257
R7228 DVSS.n2353 DVSS.n132 355.257
R7229 DVSS.n173 DVSS.n172 355.257
R7230 DVSS.n175 DVSS.n174 355.257
R7231 DVSS.n181 DVSS.n180 355.257
R7232 DVSS.n2171 DVSS.n333 355.257
R7233 DVSS.n2183 DVSS.n2182 355.257
R7234 DVSS.n2185 DVSS.n2184 355.257
R7235 DVSS.n2309 DVSS.n287 355.257
R7236 DVSS.n1989 DVSS.n405 355.257
R7237 DVSS.n2001 DVSS.n2000 355.257
R7238 DVSS.n2003 DVSS.n2002 355.257
R7239 DVSS.n2127 DVSS.n359 355.257
R7240 DVSS.n1807 DVSS.n477 355.257
R7241 DVSS.n1819 DVSS.n1818 355.257
R7242 DVSS.n1821 DVSS.n1820 355.257
R7243 DVSS.n1945 DVSS.n431 355.257
R7244 DVSS.n1000 DVSS.t116 346.384
R7245 DVSS.n1182 DVSS.t217 346.384
R7246 DVSS.n1354 DVSS.t9 346.384
R7247 DVSS.n1440 DVSS.t42 346.384
R7248 DVSS.t59 DVSS.n1570 346.384
R7249 DVSS.n1852 DVSS.t205 346.384
R7250 DVSS.n2034 DVSS.t257 346.384
R7251 DVSS.n2216 DVSS.t84 346.384
R7252 DVSS.n2388 DVSS.t255 346.384
R7253 DVSS.n2474 DVSS.t96 346.384
R7254 DVSS.t156 DVSS.n2567 346.384
R7255 DVSS.n2783 DVSS.n4 340.897
R7256 DVSS.n913 DVSS.t313 321.971
R7257 DVSS.n868 DVSS.t316 321.971
R7258 DVSS.n796 DVSS.t314 321.971
R7259 DVSS.n592 DVSS.t307 321.971
R7260 DVSS.n557 DVSS.t310 321.971
R7261 DVSS.n1603 DVSS.t309 321.971
R7262 DVSS.n448 DVSS.t312 321.971
R7263 DVSS.n376 DVSS.t311 321.971
R7264 DVSS.n304 DVSS.t308 321.971
R7265 DVSS.n100 DVSS.t315 321.971
R7266 DVSS.n65 DVSS.t317 321.971
R7267 DVSS.n1080 DVSS.t120 318.252
R7268 DVSS.n1262 DVSS.t219 318.252
R7269 DVSS.n670 DVSS.t11 318.252
R7270 DVSS.t46 DVSS.n1654 318.252
R7271 DVSS.n1753 DVSS.t61 318.252
R7272 DVSS.n2746 DVSS.t162 318.252
R7273 DVSS.t100 DVSS.n2647 318.252
R7274 DVSS.n178 DVSS.t247 318.252
R7275 DVSS.n2296 DVSS.t78 318.252
R7276 DVSS.n2114 DVSS.t267 318.252
R7277 DVSS.n1932 DVSS.t207 318.252
R7278 DVSS.t235 DVSS.n1107 317.808
R7279 DVSS.t106 DVSS.n1289 317.808
R7280 DVSS.n683 DVSS.t154 317.808
R7281 DVSS.n1696 DVSS.t188 317.808
R7282 DVSS.n2689 DVSS.t152 317.808
R7283 DVSS.n191 DVSS.t305 317.808
R7284 DVSS.t74 DVSS.n2323 317.808
R7285 DVSS.t52 DVSS.n2141 317.808
R7286 DVSS.t194 DVSS.n1959 317.808
R7287 DVSS.n1779 DVSS.t243 317.808
R7288 DVSS.t114 DVSS.n965 303.449
R7289 DVSS.t225 DVSS.n1147 303.449
R7290 DVSS.t17 DVSS.n663 303.449
R7291 DVSS.t38 DVSS.n699 303.449
R7292 DVSS.t67 DVSS.n1725 303.449
R7293 DVSS.t166 DVSS.n2718 303.449
R7294 DVSS.t104 DVSS.n207 303.449
R7295 DVSS.t253 DVSS.n171 303.449
R7296 DVSS.t82 DVSS.n2181 303.449
R7297 DVSS.t263 DVSS.n1999 303.449
R7298 DVSS.t203 DVSS.n1817 303.449
R7299 DVSS.n955 DVSS.n954 296.048
R7300 DVSS.n934 DVSS.t297 281.846
R7301 DVSS.n1057 DVSS.t282 281.846
R7302 DVSS.n1239 DVSS.t288 281.846
R7303 DVSS.n593 DVSS.t273 281.846
R7304 DVSS.n1505 DVSS.t300 281.846
R7305 DVSS.n1604 DVSS.t303 281.846
R7306 DVSS.n1909 DVSS.t291 281.846
R7307 DVSS.n2091 DVSS.t294 281.846
R7308 DVSS.n2273 DVSS.t276 281.846
R7309 DVSS.n101 DVSS.t285 281.846
R7310 DVSS.n2539 DVSS.t279 281.846
R7311 DVSS.n954 DVSS.t296 281.312
R7312 DVSS.n965 DVSS.t122 273.844
R7313 DVSS.n1147 DVSS.t223 273.844
R7314 DVSS.n663 DVSS.t13 273.844
R7315 DVSS.n699 DVSS.t44 273.844
R7316 DVSS.n1725 DVSS.t65 273.844
R7317 DVSS.n2718 DVSS.t160 273.844
R7318 DVSS.n207 DVSS.t94 273.844
R7319 DVSS.n171 DVSS.t245 273.844
R7320 DVSS.n2181 DVSS.t76 273.844
R7321 DVSS.n1999 DVSS.t261 273.844
R7322 DVSS.n1817 DVSS.t209 273.844
R7323 DVSS.n987 DVSS.n986 266.442
R7324 DVSS.n1169 DVSS.n1168 266.442
R7325 DVSS.n1340 DVSS.n1339 266.442
R7326 DVSS.n698 DVSS.n696 266.442
R7327 DVSS.n1723 DVSS.n1722 266.442
R7328 DVSS.n2716 DVSS.n2715 266.442
R7329 DVSS.n206 DVSS.n204 266.442
R7330 DVSS.n2374 DVSS.n2373 266.442
R7331 DVSS.n2203 DVSS.n2202 266.442
R7332 DVSS.n2021 DVSS.n2020 266.442
R7333 DVSS.n1839 DVSS.n1838 266.442
R7334 DVSS.n1126 DVSS.t137 263.014
R7335 DVSS.t137 DVSS.n832 263.014
R7336 DVSS.n1308 DVSS.t108 263.014
R7337 DVSS.t108 DVSS.n760 263.014
R7338 DVSS.t56 DVSS.n689 263.014
R7339 DVSS.n690 DVSS.t56 263.014
R7340 DVSS.t71 DVSS.n1708 263.014
R7341 DVSS.n1710 DVSS.t71 263.014
R7342 DVSS.t111 DVSS.n2701 263.014
R7343 DVSS.n2703 DVSS.t111 263.014
R7344 DVSS.t21 DVSS.n197 263.014
R7345 DVSS.n198 DVSS.t21 263.014
R7346 DVSS.n2342 DVSS.t202 263.014
R7347 DVSS.t202 DVSS.n268 263.014
R7348 DVSS.n2160 DVSS.t132 263.014
R7349 DVSS.t132 DVSS.n340 263.014
R7350 DVSS.n1978 DVSS.t35 263.014
R7351 DVSS.t35 DVSS.n412 263.014
R7352 DVSS.n1796 DVSS.t32 263.014
R7353 DVSS.t32 DVSS.n484 263.014
R7354 DVSS.n1077 DVSS.t281 246.553
R7355 DVSS.n1259 DVSS.t287 246.553
R7356 DVSS.n1427 DVSS.t272 246.553
R7357 DVSS.n1651 DVSS.t299 246.553
R7358 DVSS.n1584 DVSS.t302 246.553
R7359 DVSS.n1929 DVSS.t290 246.553
R7360 DVSS.n2111 DVSS.t293 246.553
R7361 DVSS.n2293 DVSS.t275 246.553
R7362 DVSS.n2461 DVSS.t284 246.553
R7363 DVSS.n2644 DVSS.t278 246.553
R7364 DVSS.n989 DVSS.n988 224.681
R7365 DVSS.n1171 DVSS.n1170 224.681
R7366 DVSS.n1342 DVSS.n1341 224.681
R7367 DVSS.n1428 DVSS.n578 224.681
R7368 DVSS.n547 DVSS.n518 224.681
R7369 DVSS.n1841 DVSS.n1840 224.681
R7370 DVSS.n2023 DVSS.n2022 224.681
R7371 DVSS.n2205 DVSS.n2204 224.681
R7372 DVSS.n2376 DVSS.n2375 224.681
R7373 DVSS.n2462 DVSS.n86 224.681
R7374 DVSS.n55 DVSS.n26 224.681
R7375 DVSS.n1080 DVSS.n1079 218.335
R7376 DVSS.n1262 DVSS.n1261 218.335
R7377 DVSS.n671 DVSS.n670 218.335
R7378 DVSS.n1654 DVSS.n1653 218.335
R7379 DVSS.n1754 DVSS.n1753 218.335
R7380 DVSS.n2747 DVSS.n2746 218.335
R7381 DVSS.n2647 DVSS.n2646 218.335
R7382 DVSS.n179 DVSS.n178 218.335
R7383 DVSS.n2296 DVSS.n2295 218.335
R7384 DVSS.n2114 DVSS.n2113 218.335
R7385 DVSS.n1932 DVSS.n1931 218.335
R7386 DVSS.n1108 DVSS.t235 208.22
R7387 DVSS.n1290 DVSS.t106 208.22
R7388 DVSS.t154 DVSS.n681 208.22
R7389 DVSS.n1681 DVSS.t188 208.22
R7390 DVSS.n2674 DVSS.t152 208.22
R7391 DVSS.t305 DVSS.n189 208.22
R7392 DVSS.n2324 DVSS.t74 208.22
R7393 DVSS.n2142 DVSS.t52 208.22
R7394 DVSS.n1960 DVSS.t194 208.22
R7395 DVSS.t243 DVSS.n1776 208.22
R7396 DVSS.n2783 DVSS.n5 200.215
R7397 DVSS.n2783 DVSS.n6 200.215
R7398 DVSS.n2783 DVSS.n7 200.215
R7399 DVSS.n2783 DVSS.n8 200.215
R7400 DVSS.n917 DVSS.n904 200.215
R7401 DVSS.n926 DVSS.n904 200.215
R7402 DVSS.n916 DVSS.n904 200.215
R7403 DVSS.n2601 DVSS.n3 200.215
R7404 DVSS.n2598 DVSS.n3 200.215
R7405 DVSS.n2588 DVSS.n3 200.215
R7406 DVSS.n2585 DVSS.n3 200.215
R7407 DVSS.n2574 DVSS.n3 200.215
R7408 DVSS.n2552 DVSS.n54 200.215
R7409 DVSS.n2550 DVSS.n54 200.215
R7410 DVSS.n2535 DVSS.n54 200.215
R7411 DVSS.n2533 DVSS.n54 200.215
R7412 DVSS.n2524 DVSS.n53 200.215
R7413 DVSS.n2522 DVSS.n53 200.215
R7414 DVSS.n2507 DVSS.n53 200.215
R7415 DVSS.n2505 DVSS.n53 200.215
R7416 DVSS.n2490 DVSS.n53 200.215
R7417 DVSS.n2460 DVSS.n2459 200.215
R7418 DVSS.n2460 DVSS.n95 200.215
R7419 DVSS.n2460 DVSS.n94 200.215
R7420 DVSS.n2460 DVSS.n93 200.215
R7421 DVSS.n2436 DVSS.n92 200.215
R7422 DVSS.n2421 DVSS.n92 200.215
R7423 DVSS.n2419 DVSS.n92 200.215
R7424 DVSS.n115 DVSS.n92 200.215
R7425 DVSS.n2404 DVSS.n92 200.215
R7426 DVSS.n2292 DVSS.n2291 200.215
R7427 DVSS.n2292 DVSS.n297 200.215
R7428 DVSS.n2292 DVSS.n296 200.215
R7429 DVSS.n2292 DVSS.n295 200.215
R7430 DVSS.n2261 DVSS.n294 200.215
R7431 DVSS.n307 DVSS.n294 200.215
R7432 DVSS.n2247 DVSS.n294 200.215
R7433 DVSS.n316 DVSS.n294 200.215
R7434 DVSS.n2232 DVSS.n294 200.215
R7435 DVSS.n2110 DVSS.n2109 200.215
R7436 DVSS.n2110 DVSS.n369 200.215
R7437 DVSS.n2110 DVSS.n368 200.215
R7438 DVSS.n2110 DVSS.n367 200.215
R7439 DVSS.n2079 DVSS.n366 200.215
R7440 DVSS.n379 DVSS.n366 200.215
R7441 DVSS.n2065 DVSS.n366 200.215
R7442 DVSS.n388 DVSS.n366 200.215
R7443 DVSS.n2050 DVSS.n366 200.215
R7444 DVSS.n1928 DVSS.n1927 200.215
R7445 DVSS.n1928 DVSS.n441 200.215
R7446 DVSS.n1928 DVSS.n440 200.215
R7447 DVSS.n1928 DVSS.n439 200.215
R7448 DVSS.n1897 DVSS.n438 200.215
R7449 DVSS.n451 DVSS.n438 200.215
R7450 DVSS.n1883 DVSS.n438 200.215
R7451 DVSS.n460 DVSS.n438 200.215
R7452 DVSS.n1868 DVSS.n438 200.215
R7453 DVSS.n1591 DVSS.n1590 200.215
R7454 DVSS.n1590 DVSS.n1589 200.215
R7455 DVSS.n1590 DVSS.n1588 200.215
R7456 DVSS.n1590 DVSS.n1586 200.215
R7457 DVSS.n1583 DVSS.n1573 200.215
R7458 DVSS.n1583 DVSS.n1576 200.215
R7459 DVSS.n1583 DVSS.n1577 200.215
R7460 DVSS.n1583 DVSS.n1580 200.215
R7461 DVSS.n1583 DVSS.n1581 200.215
R7462 DVSS.n1518 DVSS.n546 200.215
R7463 DVSS.n1516 DVSS.n546 200.215
R7464 DVSS.n1501 DVSS.n546 200.215
R7465 DVSS.n1499 DVSS.n546 200.215
R7466 DVSS.n1490 DVSS.n545 200.215
R7467 DVSS.n1488 DVSS.n545 200.215
R7468 DVSS.n1473 DVSS.n545 200.215
R7469 DVSS.n1471 DVSS.n545 200.215
R7470 DVSS.n1456 DVSS.n545 200.215
R7471 DVSS.n1426 DVSS.n1425 200.215
R7472 DVSS.n1426 DVSS.n587 200.215
R7473 DVSS.n1426 DVSS.n586 200.215
R7474 DVSS.n1426 DVSS.n585 200.215
R7475 DVSS.n1402 DVSS.n584 200.215
R7476 DVSS.n1387 DVSS.n584 200.215
R7477 DVSS.n1385 DVSS.n584 200.215
R7478 DVSS.n607 DVSS.n584 200.215
R7479 DVSS.n1370 DVSS.n584 200.215
R7480 DVSS.n1258 DVSS.n1257 200.215
R7481 DVSS.n1258 DVSS.n789 200.215
R7482 DVSS.n1258 DVSS.n788 200.215
R7483 DVSS.n1258 DVSS.n787 200.215
R7484 DVSS.n1227 DVSS.n786 200.215
R7485 DVSS.n799 DVSS.n786 200.215
R7486 DVSS.n1213 DVSS.n786 200.215
R7487 DVSS.n808 DVSS.n786 200.215
R7488 DVSS.n1198 DVSS.n786 200.215
R7489 DVSS.n1076 DVSS.n1075 200.215
R7490 DVSS.n1076 DVSS.n861 200.215
R7491 DVSS.n1076 DVSS.n860 200.215
R7492 DVSS.n1076 DVSS.n859 200.215
R7493 DVSS.n1045 DVSS.n858 200.215
R7494 DVSS.n871 DVSS.n858 200.215
R7495 DVSS.n1031 DVSS.n858 200.215
R7496 DVSS.n880 DVSS.n858 200.215
R7497 DVSS.n1016 DVSS.n858 200.215
R7498 DVSS.n953 DVSS.n952 200.215
R7499 DVSS.n953 DVSS.n906 200.215
R7500 DVSS.n953 DVSS.n905 200.215
R7501 DVSS.n969 DVSS.t118 185.03
R7502 DVSS.n1151 DVSS.t215 185.03
R7503 DVSS.n666 DVSS.t7 185.03
R7504 DVSS.t36 DVSS.n543 185.03
R7505 DVSS.t57 DVSS.n507 185.03
R7506 DVSS.t164 DVSS.n15 185.03
R7507 DVSS.t102 DVSS.n51 185.03
R7508 DVSS.n174 DVSS.t251 185.03
R7509 DVSS.n2185 DVSS.t80 185.03
R7510 DVSS.n2003 DVSS.t259 185.03
R7511 DVSS.n1821 DVSS.t213 185.03
R7512 DVSS.n928 DVSS.n916 184.572
R7513 DVSS.n926 DVSS.n925 184.572
R7514 DVSS.n917 DVSS.n903 184.572
R7515 DVSS.n2753 DVSS.n8 184.572
R7516 DVSS.n2756 DVSS.n7 184.572
R7517 DVSS.n2758 DVSS.n6 184.572
R7518 DVSS.n2759 DVSS.n5 184.572
R7519 DVSS.n2757 DVSS.n6 184.572
R7520 DVSS.n2754 DVSS.n7 184.572
R7521 DVSS.n10 DVSS.n8 184.572
R7522 DVSS.n918 DVSS.n917 184.572
R7523 DVSS.n927 DVSS.n926 184.572
R7524 DVSS.n911 DVSS.n905 184.572
R7525 DVSS.n944 DVSS.n906 184.572
R7526 DVSS.n952 DVSS.n951 184.572
R7527 DVSS.n1018 DVSS.n1016 184.572
R7528 DVSS.n1029 DVSS.n880 184.572
R7529 DVSS.n1033 DVSS.n1031 184.572
R7530 DVSS.n1043 DVSS.n871 184.572
R7531 DVSS.n1047 DVSS.n1045 184.572
R7532 DVSS.n1053 DVSS.n859 184.572
R7533 DVSS.n866 DVSS.n860 184.572
R7534 DVSS.n1067 DVSS.n861 184.572
R7535 DVSS.n1075 DVSS.n1074 184.572
R7536 DVSS.n1200 DVSS.n1198 184.572
R7537 DVSS.n1211 DVSS.n808 184.572
R7538 DVSS.n1215 DVSS.n1213 184.572
R7539 DVSS.n1225 DVSS.n799 184.572
R7540 DVSS.n1229 DVSS.n1227 184.572
R7541 DVSS.n1235 DVSS.n787 184.572
R7542 DVSS.n794 DVSS.n788 184.572
R7543 DVSS.n1249 DVSS.n789 184.572
R7544 DVSS.n1257 DVSS.n1256 184.572
R7545 DVSS.n1372 DVSS.n1370 184.572
R7546 DVSS.n1383 DVSS.n607 184.572
R7547 DVSS.n1386 DVSS.n1385 184.572
R7548 DVSS.n1387 DVSS.n599 184.572
R7549 DVSS.n1403 DVSS.n1402 184.572
R7550 DVSS.n596 DVSS.n585 184.572
R7551 DVSS.n1410 DVSS.n586 184.572
R7552 DVSS.n588 DVSS.n587 184.572
R7553 DVSS.n1425 DVSS.n582 184.572
R7554 DVSS.n1456 DVSS.n568 184.572
R7555 DVSS.n1472 DVSS.n1471 184.572
R7556 DVSS.n1473 DVSS.n562 184.572
R7557 DVSS.n1489 DVSS.n1488 184.572
R7558 DVSS.n1490 DVSS.n559 184.572
R7559 DVSS.n1500 DVSS.n1499 184.572
R7560 DVSS.n1501 DVSS.n553 184.572
R7561 DVSS.n1517 DVSS.n1516 184.572
R7562 DVSS.n1518 DVSS.n548 184.572
R7563 DVSS.n1581 DVSS.n1533 184.572
R7564 DVSS.n1580 DVSS.n1579 184.572
R7565 DVSS.n1577 DVSS.n1543 184.572
R7566 DVSS.n1576 DVSS.n1575 184.572
R7567 DVSS.n1573 DVSS.n1552 184.572
R7568 DVSS.n1586 DVSS.n1554 184.572
R7569 DVSS.n1588 DVSS.n1587 184.572
R7570 DVSS.n1589 DVSS.n1562 184.572
R7571 DVSS.n1592 DVSS.n1591 184.572
R7572 DVSS.n1870 DVSS.n1868 184.572
R7573 DVSS.n1881 DVSS.n460 184.572
R7574 DVSS.n1885 DVSS.n1883 184.572
R7575 DVSS.n1895 DVSS.n451 184.572
R7576 DVSS.n1899 DVSS.n1897 184.572
R7577 DVSS.n1905 DVSS.n439 184.572
R7578 DVSS.n446 DVSS.n440 184.572
R7579 DVSS.n1919 DVSS.n441 184.572
R7580 DVSS.n1927 DVSS.n1926 184.572
R7581 DVSS.n2052 DVSS.n2050 184.572
R7582 DVSS.n2063 DVSS.n388 184.572
R7583 DVSS.n2067 DVSS.n2065 184.572
R7584 DVSS.n2077 DVSS.n379 184.572
R7585 DVSS.n2081 DVSS.n2079 184.572
R7586 DVSS.n2087 DVSS.n367 184.572
R7587 DVSS.n374 DVSS.n368 184.572
R7588 DVSS.n2101 DVSS.n369 184.572
R7589 DVSS.n2109 DVSS.n2108 184.572
R7590 DVSS.n2234 DVSS.n2232 184.572
R7591 DVSS.n2245 DVSS.n316 184.572
R7592 DVSS.n2249 DVSS.n2247 184.572
R7593 DVSS.n2259 DVSS.n307 184.572
R7594 DVSS.n2263 DVSS.n2261 184.572
R7595 DVSS.n2269 DVSS.n295 184.572
R7596 DVSS.n302 DVSS.n296 184.572
R7597 DVSS.n2283 DVSS.n297 184.572
R7598 DVSS.n2291 DVSS.n2290 184.572
R7599 DVSS.n2406 DVSS.n2404 184.572
R7600 DVSS.n2417 DVSS.n115 184.572
R7601 DVSS.n2420 DVSS.n2419 184.572
R7602 DVSS.n2421 DVSS.n107 184.572
R7603 DVSS.n2437 DVSS.n2436 184.572
R7604 DVSS.n104 DVSS.n93 184.572
R7605 DVSS.n2444 DVSS.n94 184.572
R7606 DVSS.n96 DVSS.n95 184.572
R7607 DVSS.n2459 DVSS.n90 184.572
R7608 DVSS.n2490 DVSS.n76 184.572
R7609 DVSS.n2506 DVSS.n2505 184.572
R7610 DVSS.n2507 DVSS.n70 184.572
R7611 DVSS.n2523 DVSS.n2522 184.572
R7612 DVSS.n2524 DVSS.n67 184.572
R7613 DVSS.n2534 DVSS.n2533 184.572
R7614 DVSS.n2535 DVSS.n61 184.572
R7615 DVSS.n2551 DVSS.n2550 184.572
R7616 DVSS.n2552 DVSS.n56 184.572
R7617 DVSS.n2575 DVSS.n2574 184.572
R7618 DVSS.n2586 DVSS.n2585 184.572
R7619 DVSS.n2589 DVSS.n2588 184.572
R7620 DVSS.n2599 DVSS.n2598 184.572
R7621 DVSS.n2602 DVSS.n2601 184.572
R7622 DVSS.n2785 DVSS.n1 184.572
R7623 DVSS.n2601 DVSS.n2600 184.572
R7624 DVSS.n2598 DVSS.n2597 184.572
R7625 DVSS.n2588 DVSS.n2587 184.572
R7626 DVSS.n2585 DVSS.n2584 184.572
R7627 DVSS.n2574 DVSS.n2573 184.572
R7628 DVSS.n2553 DVSS.n2552 184.572
R7629 DVSS.n2550 DVSS.n2549 184.572
R7630 DVSS.n2536 DVSS.n2535 184.572
R7631 DVSS.n2533 DVSS.n2532 184.572
R7632 DVSS.n2525 DVSS.n2524 184.572
R7633 DVSS.n2522 DVSS.n2521 184.572
R7634 DVSS.n2508 DVSS.n2507 184.572
R7635 DVSS.n2505 DVSS.n2504 184.572
R7636 DVSS.n2491 DVSS.n2490 184.572
R7637 DVSS.n2459 DVSS.n2458 184.572
R7638 DVSS.n2445 DVSS.n95 184.572
R7639 DVSS.n105 DVSS.n94 184.572
R7640 DVSS.n2438 DVSS.n93 184.572
R7641 DVSS.n2436 DVSS.n2435 184.572
R7642 DVSS.n2422 DVSS.n2421 184.572
R7643 DVSS.n2419 DVSS.n2418 184.572
R7644 DVSS.n2405 DVSS.n115 184.572
R7645 DVSS.n2404 DVSS.n2403 184.572
R7646 DVSS.n2291 DVSS.n298 184.572
R7647 DVSS.n303 DVSS.n297 184.572
R7648 DVSS.n2270 DVSS.n296 184.572
R7649 DVSS.n2262 DVSS.n295 184.572
R7650 DVSS.n2261 DVSS.n2260 184.572
R7651 DVSS.n2248 DVSS.n307 184.572
R7652 DVSS.n2247 DVSS.n2246 184.572
R7653 DVSS.n2233 DVSS.n316 184.572
R7654 DVSS.n2232 DVSS.n2231 184.572
R7655 DVSS.n2109 DVSS.n370 184.572
R7656 DVSS.n375 DVSS.n369 184.572
R7657 DVSS.n2088 DVSS.n368 184.572
R7658 DVSS.n2080 DVSS.n367 184.572
R7659 DVSS.n2079 DVSS.n2078 184.572
R7660 DVSS.n2066 DVSS.n379 184.572
R7661 DVSS.n2065 DVSS.n2064 184.572
R7662 DVSS.n2051 DVSS.n388 184.572
R7663 DVSS.n2050 DVSS.n2049 184.572
R7664 DVSS.n1927 DVSS.n442 184.572
R7665 DVSS.n447 DVSS.n441 184.572
R7666 DVSS.n1906 DVSS.n440 184.572
R7667 DVSS.n1898 DVSS.n439 184.572
R7668 DVSS.n1897 DVSS.n1896 184.572
R7669 DVSS.n1884 DVSS.n451 184.572
R7670 DVSS.n1883 DVSS.n1882 184.572
R7671 DVSS.n1869 DVSS.n460 184.572
R7672 DVSS.n1868 DVSS.n1867 184.572
R7673 DVSS.n1591 DVSS.n1565 184.572
R7674 DVSS.n1589 DVSS.n1561 184.572
R7675 DVSS.n1588 DVSS.n1555 184.572
R7676 DVSS.n1586 DVSS.n1585 184.572
R7677 DVSS.n1573 DVSS.n1551 184.572
R7678 DVSS.n1576 DVSS.n1574 184.572
R7679 DVSS.n1577 DVSS.n1542 184.572
R7680 DVSS.n1580 DVSS.n1578 184.572
R7681 DVSS.n1581 DVSS.n1532 184.572
R7682 DVSS.n1519 DVSS.n1518 184.572
R7683 DVSS.n1516 DVSS.n1515 184.572
R7684 DVSS.n1502 DVSS.n1501 184.572
R7685 DVSS.n1499 DVSS.n1498 184.572
R7686 DVSS.n1491 DVSS.n1490 184.572
R7687 DVSS.n1488 DVSS.n1487 184.572
R7688 DVSS.n1474 DVSS.n1473 184.572
R7689 DVSS.n1471 DVSS.n1470 184.572
R7690 DVSS.n1457 DVSS.n1456 184.572
R7691 DVSS.n1425 DVSS.n1424 184.572
R7692 DVSS.n1411 DVSS.n587 184.572
R7693 DVSS.n597 DVSS.n586 184.572
R7694 DVSS.n1404 DVSS.n585 184.572
R7695 DVSS.n1402 DVSS.n1401 184.572
R7696 DVSS.n1388 DVSS.n1387 184.572
R7697 DVSS.n1385 DVSS.n1384 184.572
R7698 DVSS.n1371 DVSS.n607 184.572
R7699 DVSS.n1370 DVSS.n1369 184.572
R7700 DVSS.n1257 DVSS.n790 184.572
R7701 DVSS.n795 DVSS.n789 184.572
R7702 DVSS.n1236 DVSS.n788 184.572
R7703 DVSS.n1228 DVSS.n787 184.572
R7704 DVSS.n1227 DVSS.n1226 184.572
R7705 DVSS.n1214 DVSS.n799 184.572
R7706 DVSS.n1213 DVSS.n1212 184.572
R7707 DVSS.n1199 DVSS.n808 184.572
R7708 DVSS.n1198 DVSS.n1197 184.572
R7709 DVSS.n1075 DVSS.n862 184.572
R7710 DVSS.n867 DVSS.n861 184.572
R7711 DVSS.n1054 DVSS.n860 184.572
R7712 DVSS.n1046 DVSS.n859 184.572
R7713 DVSS.n1045 DVSS.n1044 184.572
R7714 DVSS.n1032 DVSS.n871 184.572
R7715 DVSS.n1031 DVSS.n1030 184.572
R7716 DVSS.n1017 DVSS.n880 184.572
R7717 DVSS.n1016 DVSS.n1015 184.572
R7718 DVSS.n952 DVSS.n907 184.572
R7719 DVSS.n912 DVSS.n906 184.572
R7720 DVSS.n954 DVSS.n904 173.115
R7721 DVSS.t118 DVSS.n967 170.227
R7722 DVSS.t215 DVSS.n1149 170.227
R7723 DVSS.t7 DVSS.n665 170.227
R7724 DVSS.n701 DVSS.t36 170.227
R7725 DVSS.n1727 DVSS.t57 170.227
R7726 DVSS.n2720 DVSS.t164 170.227
R7727 DVSS.n209 DVSS.t102 170.227
R7728 DVSS.t251 DVSS.n173 170.227
R7729 DVSS.t80 DVSS.n2183 170.227
R7730 DVSS.t259 DVSS.n2001 170.227
R7731 DVSS.t213 DVSS.n1819 170.227
R7732 DVSS.n1024 DVSS 161.882
R7733 DVSS.n1206 DVSS 161.882
R7734 DVSS.n1378 DVSS 161.882
R7735 DVSS.n1464 DVSS 161.882
R7736 DVSS.n1625 DVSS 161.882
R7737 DVSS.n1876 DVSS 161.882
R7738 DVSS.n2058 DVSS 161.882
R7739 DVSS.n2240 DVSS 161.882
R7740 DVSS.n2412 DVSS 161.882
R7741 DVSS.n2498 DVSS 161.882
R7742 DVSS.n2618 DVSS 161.882
R7743 DVSS.n1778 DVSS.n1777 131.507
R7744 DVSS.n939 DVSS.t298 128.196
R7745 DVSS.n1062 DVSS.t283 128.196
R7746 DVSS.n1244 DVSS.t289 128.196
R7747 DVSS.n1418 DVSS.t274 128.196
R7748 DVSS.n1511 DVSS.t301 128.196
R7749 DVSS.n1559 DVSS.t304 128.196
R7750 DVSS.n1914 DVSS.t292 128.196
R7751 DVSS.n2096 DVSS.t295 128.196
R7752 DVSS.n2278 DVSS.t277 128.196
R7753 DVSS.n2452 DVSS.t286 128.196
R7754 DVSS.n2545 DVSS.t280 128.196
R7755 DVSS.n961 DVSS.t123 116.938
R7756 DVSS.n1143 DVSS.t224 116.938
R7757 DVSS.n1325 DVSS.t14 116.938
R7758 DVSS.n716 DVSS.t45 116.938
R7759 DVSS.n1742 DVSS.t66 116.938
R7760 DVSS.n1813 DVSS.t210 116.938
R7761 DVSS.n1995 DVSS.t262 116.938
R7762 DVSS.n2177 DVSS.t77 116.938
R7763 DVSS.n2359 DVSS.t246 116.938
R7764 DVSS.n224 DVSS.t95 116.938
R7765 DVSS.n2735 DVSS.t161 116.938
R7766 DVSS DVSS.n887 113.317
R7767 DVSS DVSS.n815 113.317
R7768 DVSS DVSS.n614 113.317
R7769 DVSS DVSS.n574 113.317
R7770 DVSS DVSS.n1527 113.317
R7771 DVSS DVSS.n467 113.317
R7772 DVSS DVSS.n395 113.317
R7773 DVSS DVSS.n323 113.317
R7774 DVSS DVSS.n122 113.317
R7775 DVSS DVSS.n82 113.317
R7776 DVSS DVSS.n2561 113.317
R7777 DVSS.n883 DVSS.t173 105.028
R7778 DVSS.n811 DVSS.t199 105.028
R7779 DVSS.n610 DVSS.t148 105.028
R7780 DVSS.n570 DVSS.t233 105.028
R7781 DVSS.n1536 DVSS.t180 105.028
R7782 DVSS.n463 DVSS.t240 105.028
R7783 DVSS.n391 DVSS.t184 105.028
R7784 DVSS.n319 DVSS.t140 105.028
R7785 DVSS.n118 DVSS.t129 105.028
R7786 DVSS.n78 DVSS.t90 105.028
R7787 DVSS.n2578 DVSS.t24 105.028
R7788 DVSS.t124 DVSS.n851 96.2158
R7789 DVSS.t221 DVSS.n779 96.2158
R7790 DVSS.n672 DVSS.t15 96.2158
R7791 DVSS.n1668 DVSS.t40 96.2158
R7792 DVSS.n1755 DVSS.t63 96.2158
R7793 DVSS.n2748 DVSS.t158 96.2158
R7794 DVSS.n2661 DVSS.t98 96.2158
R7795 DVSS.n180 DVSS.t249 96.2158
R7796 DVSS.t86 DVSS.n287 96.2158
R7797 DVSS.t265 DVSS.n359 96.2158
R7798 DVSS.t211 DVSS.n431 96.2158
R7799 DVSS.n842 DVSS.n841 90.0716
R7800 DVSS.n770 DVSS.n769 90.0716
R7801 DVSS.n738 DVSS.n737 90.0716
R7802 DVSS.n1690 DVSS.n1689 90.0716
R7803 DVSS.n494 DVSS.n493 90.0716
R7804 DVSS.n422 DVSS.n421 90.0716
R7805 DVSS.n350 DVSS.n349 90.0716
R7806 DVSS.n278 DVSS.n277 90.0716
R7807 DVSS.n246 DVSS.n245 90.0716
R7808 DVSS.n2683 DVSS.n2682 90.0716
R7809 DVSS.n2767 DVSS.n2766 90.0716
R7810 DVSS.n987 DVSS.n897 88.8146
R7811 DVSS.n1169 DVSS.n825 88.8146
R7812 DVSS.n1340 DVSS.n624 88.8146
R7813 DVSS.n696 DVSS.n695 88.8146
R7814 DVSS.n1722 DVSS.n1721 88.8146
R7815 DVSS.n2715 DVSS.n2714 88.8146
R7816 DVSS.n204 DVSS.n203 88.8146
R7817 DVSS.n2374 DVSS.n132 88.8146
R7818 DVSS.n2203 DVSS.n333 88.8146
R7819 DVSS.n2021 DVSS.n405 88.8146
R7820 DVSS.n1839 DVSS.n477 88.8146
R7821 DVSS.n986 DVSS.t122 81.4135
R7822 DVSS.n1168 DVSS.t223 81.4135
R7823 DVSS.n1339 DVSS.t13 81.4135
R7824 DVSS.t44 DVSS.n698 81.4135
R7825 DVSS.t65 DVSS.n1723 81.4135
R7826 DVSS.t160 DVSS.n2716 81.4135
R7827 DVSS.t94 DVSS.n206 81.4135
R7828 DVSS.n2373 DVSS.t245 81.4135
R7829 DVSS.n2202 DVSS.t76 81.4135
R7830 DVSS.n2020 DVSS.t261 81.4135
R7831 DVSS.n1838 DVSS.t209 81.4135
R7832 DVSS.n1086 DVSS.n854 76.7239
R7833 DVSS.n961 DVSS.n854 76.7239
R7834 DVSS.n1268 DVSS.n782 76.7239
R7835 DVSS.n1143 DVSS.n782 76.7239
R7836 DVSS.n1326 DVSS.n756 76.7239
R7837 DVSS.n1326 DVSS.n1325 76.7239
R7838 DVSS.n1662 DVSS.n540 76.7239
R7839 DVSS.n716 DVSS.n540 76.7239
R7840 DVSS.n1747 DVSS.n1743 76.7239
R7841 DVSS.n1743 DVSS.n1742 76.7239
R7842 DVSS.n1938 DVSS.n434 76.7239
R7843 DVSS.n1813 DVSS.n434 76.7239
R7844 DVSS.n2120 DVSS.n362 76.7239
R7845 DVSS.n1995 DVSS.n362 76.7239
R7846 DVSS.n2302 DVSS.n290 76.7239
R7847 DVSS.n2177 DVSS.n290 76.7239
R7848 DVSS.n2360 DVSS.n264 76.7239
R7849 DVSS.n2360 DVSS.n2359 76.7239
R7850 DVSS.n2655 DVSS.n48 76.7239
R7851 DVSS.n224 DVSS.n48 76.7239
R7852 DVSS.n2740 DVSS.n2736 76.7239
R7853 DVSS.n2736 DVSS.n2735 76.7239
R7854 DVSS.n1038 DVSS 73.0358
R7855 DVSS.n1024 DVSS 73.0358
R7856 DVSS.n1220 DVSS 73.0358
R7857 DVSS.n1206 DVSS 73.0358
R7858 DVSS.n1395 DVSS 73.0358
R7859 DVSS.n1378 DVSS 73.0358
R7860 DVSS.n1480 DVSS 73.0358
R7861 DVSS.n1464 DVSS 73.0358
R7862 DVSS.n1548 DVSS 73.0358
R7863 DVSS DVSS.n1625 73.0358
R7864 DVSS.n1890 DVSS 73.0358
R7865 DVSS.n1876 DVSS 73.0358
R7866 DVSS.n2072 DVSS 73.0358
R7867 DVSS.n2058 DVSS 73.0358
R7868 DVSS.n2254 DVSS 73.0358
R7869 DVSS.n2240 DVSS 73.0358
R7870 DVSS.n2429 DVSS 73.0358
R7871 DVSS.n2412 DVSS 73.0358
R7872 DVSS.n2514 DVSS 73.0358
R7873 DVSS.n2498 DVSS 73.0358
R7874 DVSS.n2594 DVSS 73.0358
R7875 DVSS DVSS.n2618 73.0358
R7876 DVSS.n1106 DVSS.t112 60.2745
R7877 DVSS.n1288 DVSS.t190 60.2745
R7878 DVSS.t28 DVSS.n684 60.2745
R7879 DVSS.t30 DVSS.n1697 60.2745
R7880 DVSS.t72 DVSS.n2690 60.2745
R7881 DVSS.t227 DVSS.n192 60.2745
R7882 DVSS.n2322 DVSS.t192 60.2745
R7883 DVSS.n2140 DVSS.t4 60.2745
R7884 DVSS.n1958 DVSS.t144 60.2745
R7885 DVSS.n1777 DVSS.t109 60.2745
R7886 DVSS.n1039 DVSS.n874 57.0829
R7887 DVSS.n1221 DVSS.n802 57.0829
R7888 DVSS.n1396 DVSS.n601 57.0829
R7889 DVSS.n1483 DVSS.n564 57.0829
R7890 DVSS.n1616 DVSS.n1545 57.0829
R7891 DVSS.n1891 DVSS.n454 57.0829
R7892 DVSS.n2073 DVSS.n382 57.0829
R7893 DVSS.n2255 DVSS.n310 57.0829
R7894 DVSS.n2430 DVSS.n109 57.0829
R7895 DVSS.n2517 DVSS.n72 57.0829
R7896 DVSS.n2609 DVSS.n2591 57.0829
R7897 DVSS.n1086 DVSS.n1085 57.0817
R7898 DVSS.n976 DVSS.n975 57.0817
R7899 DVSS.n1268 DVSS.n1267 57.0817
R7900 DVSS.n1158 DVSS.n1157 57.0817
R7901 DVSS.n756 DVSS.n633 57.0817
R7902 DVSS.n1329 DVSS.n1328 57.0817
R7903 DVSS.n1662 DVSS.n1661 57.0817
R7904 DVSS.n708 DVSS.n704 57.0817
R7905 DVSS.n1747 DVSS.n1744 57.0817
R7906 DVSS.n511 DVSS.n510 57.0817
R7907 DVSS.n1938 DVSS.n1937 57.0817
R7908 DVSS.n1828 DVSS.n1827 57.0817
R7909 DVSS.n2120 DVSS.n2119 57.0817
R7910 DVSS.n2010 DVSS.n2009 57.0817
R7911 DVSS.n2302 DVSS.n2301 57.0817
R7912 DVSS.n2192 DVSS.n2191 57.0817
R7913 DVSS.n264 DVSS.n141 57.0817
R7914 DVSS.n2363 DVSS.n2362 57.0817
R7915 DVSS.n2655 DVSS.n2654 57.0817
R7916 DVSS.n216 DVSS.n212 57.0817
R7917 DVSS.n2740 DVSS.n2737 57.0817
R7918 DVSS.n19 DVSS.n18 57.0817
R7919 DVSS.n1078 DVSS.n1077 52.3335
R7920 DVSS.n1260 DVSS.n1259 52.3335
R7921 DVSS.n1427 DVSS.n583 52.3335
R7922 DVSS.n1652 DVSS.n1651 52.3335
R7923 DVSS.n1584 DVSS.n1572 52.3335
R7924 DVSS.n1930 DVSS.n1929 52.3335
R7925 DVSS.n2112 DVSS.n2111 52.3335
R7926 DVSS.n2294 DVSS.n2293 52.3335
R7927 DVSS.n2461 DVSS.n91 52.3335
R7928 DVSS.n2645 DVSS.n2644 52.3335
R7929 DVSS.n2784 DVSS.n2 52.3335
R7930 DVSS.n966 DVSS.t114 51.8087
R7931 DVSS.n1148 DVSS.t225 51.8087
R7932 DVSS.n664 DVSS.t17 51.8087
R7933 DVSS.n700 DVSS.t38 51.8087
R7934 DVSS.n1726 DVSS.t67 51.8087
R7935 DVSS.n2719 DVSS.t166 51.8087
R7936 DVSS.n208 DVSS.t104 51.8087
R7937 DVSS.n172 DVSS.t253 51.8087
R7938 DVSS.n2182 DVSS.t82 51.8087
R7939 DVSS.n2000 DVSS.t263 51.8087
R7940 DVSS.n1818 DVSS.t203 51.8087
R7941 DVSS.n877 DVSS.n876 46.2505
R7942 DVSS.n805 DVSS.n804 46.2505
R7943 DVSS.n605 DVSS.n604 46.2505
R7944 DVSS.n566 DVSS.n565 46.2505
R7945 DVSS.n1538 DVSS.n1537 46.2505
R7946 DVSS.n457 DVSS.n456 46.2505
R7947 DVSS.n385 DVSS.n384 46.2505
R7948 DVSS.n313 DVSS.n312 46.2505
R7949 DVSS.n113 DVSS.n112 46.2505
R7950 DVSS.n74 DVSS.n73 46.2505
R7951 DVSS.n2580 DVSS.n2579 46.2505
R7952 DVSS.n1038 DVSS 44.424
R7953 DVSS.n1220 DVSS 44.424
R7954 DVSS.n1395 DVSS 44.424
R7955 DVSS.n1480 DVSS 44.424
R7956 DVSS.n1548 DVSS 44.424
R7957 DVSS.n1890 DVSS 44.424
R7958 DVSS.n2072 DVSS 44.424
R7959 DVSS.n2254 DVSS 44.424
R7960 DVSS.n2429 DVSS 44.424
R7961 DVSS.n2514 DVSS 44.424
R7962 DVSS.n2594 DVSS 44.424
R7963 DVSS.n1079 DVSS.t124 40.707
R7964 DVSS.n1261 DVSS.t221 40.707
R7965 DVSS.t15 DVSS.n671 40.707
R7966 DVSS.n1653 DVSS.t40 40.707
R7967 DVSS.t63 DVSS.n1754 40.707
R7968 DVSS.t158 DVSS.n2747 40.707
R7969 DVSS.n2646 DVSS.t98 40.707
R7970 DVSS.t249 DVSS.n179 40.707
R7971 DVSS.n2295 DVSS.t86 40.707
R7972 DVSS.n2113 DVSS.t265 40.707
R7973 DVSS.n1931 DVSS.t211 40.707
R7974 DVSS.n968 DVSS.t120 37.0064
R7975 DVSS.n1150 DVSS.t219 37.0064
R7976 DVSS.n667 DVSS.t11 37.0064
R7977 DVSS.n1655 DVSS.t46 37.0064
R7978 DVSS.t61 DVSS.n1752 37.0064
R7979 DVSS.t162 DVSS.n2745 37.0064
R7980 DVSS.n2648 DVSS.t100 37.0064
R7981 DVSS.n175 DVSS.t247 37.0064
R7982 DVSS.n2184 DVSS.t78 37.0064
R7983 DVSS.n2002 DVSS.t267 37.0064
R7984 DVSS.n1820 DVSS.t207 37.0064
R7985 DVSS.n932 DVSS.n910 36.1417
R7986 DVSS.n943 DVSS.n910 36.1417
R7987 DVSS.n945 DVSS.n943 36.1417
R7988 DVSS.n945 DVSS.n908 36.1417
R7989 DVSS.n950 DVSS.n908 36.1417
R7990 DVSS.n950 DVSS.n894 36.1417
R7991 DVSS.n991 DVSS.n894 36.1417
R7992 DVSS.n991 DVSS.n893 36.1417
R7993 DVSS.n996 DVSS.n893 36.1417
R7994 DVSS.n996 DVSS.n889 36.1417
R7995 DVSS.n1002 DVSS.n889 36.1417
R7996 DVSS.n1002 DVSS.n886 36.1417
R7997 DVSS.n1013 DVSS.n886 36.1417
R7998 DVSS.n1013 DVSS.n884 36.1417
R7999 DVSS.n1019 DVSS.n884 36.1417
R8000 DVSS.n1019 DVSS.n881 36.1417
R8001 DVSS.n1028 DVSS.n881 36.1417
R8002 DVSS.n1028 DVSS.n879 36.1417
R8003 DVSS.n1034 DVSS.n879 36.1417
R8004 DVSS.n1034 DVSS.n872 36.1417
R8005 DVSS.n1042 DVSS.n872 36.1417
R8006 DVSS.n1042 DVSS.n870 36.1417
R8007 DVSS.n1048 DVSS.n870 36.1417
R8008 DVSS.n1048 DVSS.n869 36.1417
R8009 DVSS.n1052 DVSS.n869 36.1417
R8010 DVSS.n1055 DVSS.n1052 36.1417
R8011 DVSS.n1055 DVSS.n865 36.1417
R8012 DVSS.n1066 DVSS.n865 36.1417
R8013 DVSS.n1068 DVSS.n1066 36.1417
R8014 DVSS.n1068 DVSS.n863 36.1417
R8015 DVSS.n1073 DVSS.n863 36.1417
R8016 DVSS.n1073 DVSS.n822 36.1417
R8017 DVSS.n1173 DVSS.n822 36.1417
R8018 DVSS.n1173 DVSS.n821 36.1417
R8019 DVSS.n1178 DVSS.n821 36.1417
R8020 DVSS.n1178 DVSS.n817 36.1417
R8021 DVSS.n1184 DVSS.n817 36.1417
R8022 DVSS.n1184 DVSS.n814 36.1417
R8023 DVSS.n1195 DVSS.n814 36.1417
R8024 DVSS.n1195 DVSS.n812 36.1417
R8025 DVSS.n1201 DVSS.n812 36.1417
R8026 DVSS.n1201 DVSS.n809 36.1417
R8027 DVSS.n1210 DVSS.n809 36.1417
R8028 DVSS.n1210 DVSS.n807 36.1417
R8029 DVSS.n1216 DVSS.n807 36.1417
R8030 DVSS.n1216 DVSS.n800 36.1417
R8031 DVSS.n1224 DVSS.n800 36.1417
R8032 DVSS.n1224 DVSS.n798 36.1417
R8033 DVSS.n1230 DVSS.n798 36.1417
R8034 DVSS.n1230 DVSS.n797 36.1417
R8035 DVSS.n1234 DVSS.n797 36.1417
R8036 DVSS.n1237 DVSS.n1234 36.1417
R8037 DVSS.n1237 DVSS.n793 36.1417
R8038 DVSS.n1248 DVSS.n793 36.1417
R8039 DVSS.n1250 DVSS.n1248 36.1417
R8040 DVSS.n1250 DVSS.n791 36.1417
R8041 DVSS.n1255 DVSS.n791 36.1417
R8042 DVSS.n1255 DVSS.n621 36.1417
R8043 DVSS.n1344 DVSS.n621 36.1417
R8044 DVSS.n1344 DVSS.n620 36.1417
R8045 DVSS.n1349 DVSS.n620 36.1417
R8046 DVSS.n1349 DVSS.n616 36.1417
R8047 DVSS.n1356 DVSS.n616 36.1417
R8048 DVSS.n1356 DVSS.n613 36.1417
R8049 DVSS.n1367 DVSS.n613 36.1417
R8050 DVSS.n1367 DVSS.n611 36.1417
R8051 DVSS.n1373 DVSS.n611 36.1417
R8052 DVSS.n1373 DVSS.n608 36.1417
R8053 DVSS.n1382 DVSS.n608 36.1417
R8054 DVSS.n1382 DVSS.n606 36.1417
R8055 DVSS.n1391 DVSS.n606 36.1417
R8056 DVSS.n1391 DVSS.n1390 36.1417
R8057 DVSS.n1390 DVSS.n600 36.1417
R8058 DVSS.n1400 DVSS.n600 36.1417
R8059 DVSS.n1400 DVSS.n598 36.1417
R8060 DVSS.n1405 DVSS.n598 36.1417
R8061 DVSS.n1405 DVSS.n595 36.1417
R8062 DVSS.n1409 DVSS.n595 36.1417
R8063 DVSS.n1413 DVSS.n1409 36.1417
R8064 DVSS.n1413 DVSS.n1412 36.1417
R8065 DVSS.n1412 DVSS.n589 36.1417
R8066 DVSS.n1423 DVSS.n589 36.1417
R8067 DVSS.n1423 DVSS.n581 36.1417
R8068 DVSS.n1431 DVSS.n581 36.1417
R8069 DVSS.n1431 DVSS.n580 36.1417
R8070 DVSS.n1436 DVSS.n580 36.1417
R8071 DVSS.n1436 DVSS.n576 36.1417
R8072 DVSS.n1443 DVSS.n576 36.1417
R8073 DVSS.n1443 DVSS.n573 36.1417
R8074 DVSS.n1453 DVSS.n573 36.1417
R8075 DVSS.n1453 DVSS.n571 36.1417
R8076 DVSS.n1458 DVSS.n571 36.1417
R8077 DVSS.n1458 DVSS.n569 36.1417
R8078 DVSS.n1469 DVSS.n569 36.1417
R8079 DVSS.n1469 DVSS.n567 36.1417
R8080 DVSS.n1475 DVSS.n567 36.1417
R8081 DVSS.n1475 DVSS.n563 36.1417
R8082 DVSS.n1486 DVSS.n563 36.1417
R8083 DVSS.n1486 DVSS.n561 36.1417
R8084 DVSS.n1492 DVSS.n561 36.1417
R8085 DVSS.n1492 DVSS.n560 36.1417
R8086 DVSS.n1497 DVSS.n560 36.1417
R8087 DVSS.n1497 DVSS.n558 36.1417
R8088 DVSS.n1503 DVSS.n558 36.1417
R8089 DVSS.n1503 DVSS.n554 36.1417
R8090 DVSS.n1514 DVSS.n554 36.1417
R8091 DVSS.n1514 DVSS.n552 36.1417
R8092 DVSS.n1520 DVSS.n552 36.1417
R8093 DVSS.n1520 DVSS.n550 36.1417
R8094 DVSS.n1648 DVSS.n550 36.1417
R8095 DVSS.n1648 DVSS.n551 36.1417
R8096 DVSS.n1644 DVSS.n551 36.1417
R8097 DVSS.n1644 DVSS.n1643 36.1417
R8098 DVSS.n1643 DVSS.n1525 36.1417
R8099 DVSS.n1635 DVSS.n1525 36.1417
R8100 DVSS.n1635 DVSS.n1634 36.1417
R8101 DVSS.n1634 DVSS.n1530 36.1417
R8102 DVSS.n1630 DVSS.n1530 36.1417
R8103 DVSS.n1630 DVSS.n1629 36.1417
R8104 DVSS.n1629 DVSS.n1534 36.1417
R8105 DVSS.n1541 DVSS.n1534 36.1417
R8106 DVSS.n1621 DVSS.n1541 36.1417
R8107 DVSS.n1621 DVSS.n1620 36.1417
R8108 DVSS.n1620 DVSS.n1544 36.1417
R8109 DVSS.n1550 DVSS.n1544 36.1417
R8110 DVSS.n1613 DVSS.n1550 36.1417
R8111 DVSS.n1613 DVSS.n1612 36.1417
R8112 DVSS.n1612 DVSS.n1553 36.1417
R8113 DVSS.n1608 DVSS.n1553 36.1417
R8114 DVSS.n1608 DVSS.n1607 36.1417
R8115 DVSS.n1607 DVSS.n1556 36.1417
R8116 DVSS.n1598 DVSS.n1556 36.1417
R8117 DVSS.n1598 DVSS.n1597 36.1417
R8118 DVSS.n1597 DVSS.n1563 36.1417
R8119 DVSS.n1593 DVSS.n1563 36.1417
R8120 DVSS.n1593 DVSS.n474 36.1417
R8121 DVSS.n1843 DVSS.n474 36.1417
R8122 DVSS.n1843 DVSS.n473 36.1417
R8123 DVSS.n1848 DVSS.n473 36.1417
R8124 DVSS.n1848 DVSS.n469 36.1417
R8125 DVSS.n1854 DVSS.n469 36.1417
R8126 DVSS.n1854 DVSS.n466 36.1417
R8127 DVSS.n1865 DVSS.n466 36.1417
R8128 DVSS.n1865 DVSS.n464 36.1417
R8129 DVSS.n1871 DVSS.n464 36.1417
R8130 DVSS.n1871 DVSS.n461 36.1417
R8131 DVSS.n1880 DVSS.n461 36.1417
R8132 DVSS.n1880 DVSS.n459 36.1417
R8133 DVSS.n1886 DVSS.n459 36.1417
R8134 DVSS.n1886 DVSS.n452 36.1417
R8135 DVSS.n1894 DVSS.n452 36.1417
R8136 DVSS.n1894 DVSS.n450 36.1417
R8137 DVSS.n1900 DVSS.n450 36.1417
R8138 DVSS.n1900 DVSS.n449 36.1417
R8139 DVSS.n1904 DVSS.n449 36.1417
R8140 DVSS.n1907 DVSS.n1904 36.1417
R8141 DVSS.n1907 DVSS.n445 36.1417
R8142 DVSS.n1918 DVSS.n445 36.1417
R8143 DVSS.n1920 DVSS.n1918 36.1417
R8144 DVSS.n1920 DVSS.n443 36.1417
R8145 DVSS.n1925 DVSS.n443 36.1417
R8146 DVSS.n1925 DVSS.n402 36.1417
R8147 DVSS.n2025 DVSS.n402 36.1417
R8148 DVSS.n2025 DVSS.n401 36.1417
R8149 DVSS.n2030 DVSS.n401 36.1417
R8150 DVSS.n2030 DVSS.n397 36.1417
R8151 DVSS.n2036 DVSS.n397 36.1417
R8152 DVSS.n2036 DVSS.n394 36.1417
R8153 DVSS.n2047 DVSS.n394 36.1417
R8154 DVSS.n2047 DVSS.n392 36.1417
R8155 DVSS.n2053 DVSS.n392 36.1417
R8156 DVSS.n2053 DVSS.n389 36.1417
R8157 DVSS.n2062 DVSS.n389 36.1417
R8158 DVSS.n2062 DVSS.n387 36.1417
R8159 DVSS.n2068 DVSS.n387 36.1417
R8160 DVSS.n2068 DVSS.n380 36.1417
R8161 DVSS.n2076 DVSS.n380 36.1417
R8162 DVSS.n2076 DVSS.n378 36.1417
R8163 DVSS.n2082 DVSS.n378 36.1417
R8164 DVSS.n2082 DVSS.n377 36.1417
R8165 DVSS.n2086 DVSS.n377 36.1417
R8166 DVSS.n2089 DVSS.n2086 36.1417
R8167 DVSS.n2089 DVSS.n373 36.1417
R8168 DVSS.n2100 DVSS.n373 36.1417
R8169 DVSS.n2102 DVSS.n2100 36.1417
R8170 DVSS.n2102 DVSS.n371 36.1417
R8171 DVSS.n2107 DVSS.n371 36.1417
R8172 DVSS.n2107 DVSS.n330 36.1417
R8173 DVSS.n2207 DVSS.n330 36.1417
R8174 DVSS.n2207 DVSS.n329 36.1417
R8175 DVSS.n2212 DVSS.n329 36.1417
R8176 DVSS.n2212 DVSS.n325 36.1417
R8177 DVSS.n2218 DVSS.n325 36.1417
R8178 DVSS.n2218 DVSS.n322 36.1417
R8179 DVSS.n2229 DVSS.n322 36.1417
R8180 DVSS.n2229 DVSS.n320 36.1417
R8181 DVSS.n2235 DVSS.n320 36.1417
R8182 DVSS.n2235 DVSS.n317 36.1417
R8183 DVSS.n2244 DVSS.n317 36.1417
R8184 DVSS.n2244 DVSS.n315 36.1417
R8185 DVSS.n2250 DVSS.n315 36.1417
R8186 DVSS.n2250 DVSS.n308 36.1417
R8187 DVSS.n2258 DVSS.n308 36.1417
R8188 DVSS.n2258 DVSS.n306 36.1417
R8189 DVSS.n2264 DVSS.n306 36.1417
R8190 DVSS.n2264 DVSS.n305 36.1417
R8191 DVSS.n2268 DVSS.n305 36.1417
R8192 DVSS.n2271 DVSS.n2268 36.1417
R8193 DVSS.n2271 DVSS.n301 36.1417
R8194 DVSS.n2282 DVSS.n301 36.1417
R8195 DVSS.n2284 DVSS.n2282 36.1417
R8196 DVSS.n2284 DVSS.n299 36.1417
R8197 DVSS.n2289 DVSS.n299 36.1417
R8198 DVSS.n2289 DVSS.n129 36.1417
R8199 DVSS.n2378 DVSS.n129 36.1417
R8200 DVSS.n2378 DVSS.n128 36.1417
R8201 DVSS.n2383 DVSS.n128 36.1417
R8202 DVSS.n2383 DVSS.n124 36.1417
R8203 DVSS.n2390 DVSS.n124 36.1417
R8204 DVSS.n2390 DVSS.n121 36.1417
R8205 DVSS.n2401 DVSS.n121 36.1417
R8206 DVSS.n2401 DVSS.n119 36.1417
R8207 DVSS.n2407 DVSS.n119 36.1417
R8208 DVSS.n2407 DVSS.n116 36.1417
R8209 DVSS.n2416 DVSS.n116 36.1417
R8210 DVSS.n2416 DVSS.n114 36.1417
R8211 DVSS.n2425 DVSS.n114 36.1417
R8212 DVSS.n2425 DVSS.n2424 36.1417
R8213 DVSS.n2424 DVSS.n108 36.1417
R8214 DVSS.n2434 DVSS.n108 36.1417
R8215 DVSS.n2434 DVSS.n106 36.1417
R8216 DVSS.n2439 DVSS.n106 36.1417
R8217 DVSS.n2439 DVSS.n103 36.1417
R8218 DVSS.n2443 DVSS.n103 36.1417
R8219 DVSS.n2447 DVSS.n2443 36.1417
R8220 DVSS.n2447 DVSS.n2446 36.1417
R8221 DVSS.n2446 DVSS.n97 36.1417
R8222 DVSS.n2457 DVSS.n97 36.1417
R8223 DVSS.n2457 DVSS.n89 36.1417
R8224 DVSS.n2465 DVSS.n89 36.1417
R8225 DVSS.n2465 DVSS.n88 36.1417
R8226 DVSS.n2470 DVSS.n88 36.1417
R8227 DVSS.n2470 DVSS.n84 36.1417
R8228 DVSS.n2477 DVSS.n84 36.1417
R8229 DVSS.n2477 DVSS.n81 36.1417
R8230 DVSS.n2487 DVSS.n81 36.1417
R8231 DVSS.n2487 DVSS.n79 36.1417
R8232 DVSS.n2492 DVSS.n79 36.1417
R8233 DVSS.n2492 DVSS.n77 36.1417
R8234 DVSS.n2503 DVSS.n77 36.1417
R8235 DVSS.n2503 DVSS.n75 36.1417
R8236 DVSS.n2509 DVSS.n75 36.1417
R8237 DVSS.n2509 DVSS.n71 36.1417
R8238 DVSS.n2520 DVSS.n71 36.1417
R8239 DVSS.n2520 DVSS.n69 36.1417
R8240 DVSS.n2526 DVSS.n69 36.1417
R8241 DVSS.n2526 DVSS.n68 36.1417
R8242 DVSS.n2531 DVSS.n68 36.1417
R8243 DVSS.n2531 DVSS.n66 36.1417
R8244 DVSS.n2537 DVSS.n66 36.1417
R8245 DVSS.n2537 DVSS.n62 36.1417
R8246 DVSS.n2548 DVSS.n62 36.1417
R8247 DVSS.n2548 DVSS.n60 36.1417
R8248 DVSS.n2554 DVSS.n60 36.1417
R8249 DVSS.n2554 DVSS.n58 36.1417
R8250 DVSS.n2641 DVSS.n58 36.1417
R8251 DVSS.n2641 DVSS.n59 36.1417
R8252 DVSS.n2637 DVSS.n59 36.1417
R8253 DVSS.n2637 DVSS.n2636 36.1417
R8254 DVSS.n2636 DVSS.n2559 36.1417
R8255 DVSS.n2628 DVSS.n2559 36.1417
R8256 DVSS.n2628 DVSS.n2627 36.1417
R8257 DVSS.n2627 DVSS.n2570 36.1417
R8258 DVSS.n2623 DVSS.n2570 36.1417
R8259 DVSS.n2623 DVSS.n2622 36.1417
R8260 DVSS.n2622 DVSS.n2576 36.1417
R8261 DVSS.n2583 DVSS.n2576 36.1417
R8262 DVSS.n2614 DVSS.n2583 36.1417
R8263 DVSS.n2614 DVSS.n2613 36.1417
R8264 DVSS.n2613 DVSS.n2590 36.1417
R8265 DVSS.n2596 DVSS.n2590 36.1417
R8266 DVSS.n2606 DVSS.n2596 36.1417
R8267 DVSS.n2606 DVSS.n2605 36.1417
R8268 DVSS.n2605 DVSS.n0 36.1417
R8269 DVSS.n2786 DVSS.n0 36.1417
R8270 DVSS.n1006 DVSS 33.9483
R8271 DVSS.n1188 DVSS 33.9483
R8272 DVSS.n1360 DVSS 33.9483
R8273 DVSS.n1448 DVSS 33.9483
R8274 DVSS.n1639 DVSS 33.9483
R8275 DVSS.n1858 DVSS 33.9483
R8276 DVSS.n2040 DVSS 33.9483
R8277 DVSS.n2222 DVSS 33.9483
R8278 DVSS.n2394 DVSS 33.9483
R8279 DVSS.n2482 DVSS 33.9483
R8280 DVSS.n2632 DVSS 33.9483
R8281 DVSS.n841 DVSS.t236 28.1205
R8282 DVSS.n769 DVSS.t107 28.1205
R8283 DVSS.n737 DVSS.t155 28.1205
R8284 DVSS.n1689 DVSS.t189 28.1205
R8285 DVSS.n493 DVSS.t244 28.1205
R8286 DVSS.n421 DVSS.t195 28.1205
R8287 DVSS.n349 DVSS.t53 28.1205
R8288 DVSS.n277 DVSS.t75 28.1205
R8289 DVSS.n245 DVSS.t306 28.1205
R8290 DVSS.n2682 DVSS.t153 28.1205
R8291 DVSS.n2766 DVSS.t6 28.1205
R8292 DVSS.n1006 DVSS.n1005 21.8222
R8293 DVSS.n1188 DVSS.n1187 21.8222
R8294 DVSS.n1360 DVSS.n1359 21.8222
R8295 DVSS.n1448 DVSS.n1447 21.8222
R8296 DVSS.n1640 DVSS.n1639 21.8222
R8297 DVSS.n1858 DVSS.n1857 21.8222
R8298 DVSS.n2040 DVSS.n2039 21.8222
R8299 DVSS.n2222 DVSS.n2221 21.8222
R8300 DVSS.n2394 DVSS.n2393 21.8222
R8301 DVSS.n2482 DVSS.n2481 21.8222
R8302 DVSS.n2633 DVSS.n2632 21.8222
R8303 DVSS.n841 DVSS.t113 21.2805
R8304 DVSS.n769 DVSS.t191 21.2805
R8305 DVSS.n737 DVSS.t29 21.2805
R8306 DVSS.n1689 DVSS.t31 21.2805
R8307 DVSS.n493 DVSS.t110 21.2805
R8308 DVSS.n421 DVSS.t145 21.2805
R8309 DVSS.n349 DVSS.t5 21.2805
R8310 DVSS.n277 DVSS.t193 21.2805
R8311 DVSS.n245 DVSS.t228 21.2805
R8312 DVSS.n2682 DVSS.t73 21.2805
R8313 DVSS.n2766 DVSS.t3 21.2805
R8314 DVSS.n887 DVSS.t271 20.0005
R8315 DVSS.n887 DVSS.t117 20.0005
R8316 DVSS.n815 DVSS.t136 20.0005
R8317 DVSS.n815 DVSS.t218 20.0005
R8318 DVSS.n614 DVSS.t1 20.0005
R8319 DVSS.n614 DVSS.t10 20.0005
R8320 DVSS.n574 DVSS.t55 20.0005
R8321 DVSS.n574 DVSS.t43 20.0005
R8322 DVSS.n1527 DVSS.t70 20.0005
R8323 DVSS.n1527 DVSS.t60 20.0005
R8324 DVSS.n467 DVSS.t49 20.0005
R8325 DVSS.n467 DVSS.t206 20.0005
R8326 DVSS.n395 DVSS.t34 20.0005
R8327 DVSS.n395 DVSS.t258 20.0005
R8328 DVSS.n323 DVSS.t134 20.0005
R8329 DVSS.n323 DVSS.t85 20.0005
R8330 DVSS.n122 DVSS.t51 20.0005
R8331 DVSS.n122 DVSS.t256 20.0005
R8332 DVSS.n82 DVSS.t20 20.0005
R8333 DVSS.n82 DVSS.t97 20.0005
R8334 DVSS.n2561 DVSS.t169 20.0005
R8335 DVSS.n2561 DVSS.t157 20.0005
R8336 DVSS.n935 DVSS.n934 14.5464
R8337 DVSS.n1058 DVSS.n1057 14.5464
R8338 DVSS.n1240 DVSS.n1239 14.5464
R8339 DVSS.n594 DVSS.n593 14.5464
R8340 DVSS.n1506 DVSS.n1505 14.5464
R8341 DVSS.n1605 DVSS.n1604 14.5464
R8342 DVSS.n1910 DVSS.n1909 14.5464
R8343 DVSS.n2092 DVSS.n2091 14.5464
R8344 DVSS.n2274 DVSS.n2273 14.5464
R8345 DVSS.n102 DVSS.n101 14.5464
R8346 DVSS.n2540 DVSS.n2539 14.5464
R8347 DVSS.n1007 DVSS.n1006 12.5222
R8348 DVSS.n1189 DVSS.n1188 12.5222
R8349 DVSS.n1361 DVSS.n1360 12.5222
R8350 DVSS.n1449 DVSS.n1448 12.5222
R8351 DVSS.n1639 DVSS.n1526 12.5222
R8352 DVSS.n1859 DVSS.n1858 12.5222
R8353 DVSS.n2041 DVSS.n2040 12.5222
R8354 DVSS.n2223 DVSS.n2222 12.5222
R8355 DVSS.n2395 DVSS.n2394 12.5222
R8356 DVSS.n2483 DVSS.n2482 12.5222
R8357 DVSS.n2632 DVSS.n2560 12.5222
R8358 DVSS.n1085 DVSS.t121 10.6405
R8359 DVSS.n1085 DVSS.t125 10.6405
R8360 DVSS.n975 DVSS.t115 10.6405
R8361 DVSS.n975 DVSS.t119 10.6405
R8362 DVSS.n1267 DVSS.t220 10.6405
R8363 DVSS.n1267 DVSS.t222 10.6405
R8364 DVSS.n1157 DVSS.t226 10.6405
R8365 DVSS.n1157 DVSS.t216 10.6405
R8366 DVSS.n633 DVSS.t12 10.6405
R8367 DVSS.n633 DVSS.t16 10.6405
R8368 DVSS.n1328 DVSS.t18 10.6405
R8369 DVSS.n1328 DVSS.t8 10.6405
R8370 DVSS.n1661 DVSS.t47 10.6405
R8371 DVSS.n1661 DVSS.t41 10.6405
R8372 DVSS.n704 DVSS.t39 10.6405
R8373 DVSS.n704 DVSS.t37 10.6405
R8374 DVSS.n1744 DVSS.t62 10.6405
R8375 DVSS.n1744 DVSS.t64 10.6405
R8376 DVSS.n510 DVSS.t68 10.6405
R8377 DVSS.n510 DVSS.t58 10.6405
R8378 DVSS.n1937 DVSS.t208 10.6405
R8379 DVSS.n1937 DVSS.t212 10.6405
R8380 DVSS.n1827 DVSS.t204 10.6405
R8381 DVSS.n1827 DVSS.t214 10.6405
R8382 DVSS.n2119 DVSS.t268 10.6405
R8383 DVSS.n2119 DVSS.t266 10.6405
R8384 DVSS.n2009 DVSS.t264 10.6405
R8385 DVSS.n2009 DVSS.t260 10.6405
R8386 DVSS.n2301 DVSS.t79 10.6405
R8387 DVSS.n2301 DVSS.t87 10.6405
R8388 DVSS.n2191 DVSS.t83 10.6405
R8389 DVSS.n2191 DVSS.t81 10.6405
R8390 DVSS.n141 DVSS.t248 10.6405
R8391 DVSS.n141 DVSS.t250 10.6405
R8392 DVSS.n2362 DVSS.t254 10.6405
R8393 DVSS.n2362 DVSS.t252 10.6405
R8394 DVSS.n2654 DVSS.t101 10.6405
R8395 DVSS.n2654 DVSS.t99 10.6405
R8396 DVSS.n212 DVSS.t105 10.6405
R8397 DVSS.n212 DVSS.t103 10.6405
R8398 DVSS.n2737 DVSS.t163 10.6405
R8399 DVSS.n2737 DVSS.t159 10.6405
R8400 DVSS.n18 DVSS.t167 10.6405
R8401 DVSS.n18 DVSS.t165 10.6405
R8402 DVSS.n876 DVSS.t175 10.6405
R8403 DVSS.n876 DVSS.t171 10.6405
R8404 DVSS.n874 DVSS.t172 10.6405
R8405 DVSS.n874 DVSS.t174 10.6405
R8406 DVSS.n804 DVSS.t201 10.6405
R8407 DVSS.n804 DVSS.t200 10.6405
R8408 DVSS.n802 DVSS.t198 10.6405
R8409 DVSS.n802 DVSS.t197 10.6405
R8410 DVSS.n604 DVSS.t149 10.6405
R8411 DVSS.n604 DVSS.t151 10.6405
R8412 DVSS.n601 DVSS.t147 10.6405
R8413 DVSS.n601 DVSS.t150 10.6405
R8414 DVSS.n565 DVSS.t231 10.6405
R8415 DVSS.n565 DVSS.t230 10.6405
R8416 DVSS.n564 DVSS.t232 10.6405
R8417 DVSS.n564 DVSS.t234 10.6405
R8418 DVSS.n1537 DVSS.t181 10.6405
R8419 DVSS.n1537 DVSS.t177 10.6405
R8420 DVSS.n1545 DVSS.t178 10.6405
R8421 DVSS.n1545 DVSS.t179 10.6405
R8422 DVSS.n456 DVSS.t242 10.6405
R8423 DVSS.n456 DVSS.t238 10.6405
R8424 DVSS.n454 DVSS.t239 10.6405
R8425 DVSS.n454 DVSS.t241 10.6405
R8426 DVSS.n384 DVSS.t187 10.6405
R8427 DVSS.n384 DVSS.t186 10.6405
R8428 DVSS.n382 DVSS.t183 10.6405
R8429 DVSS.n382 DVSS.t185 10.6405
R8430 DVSS.n312 DVSS.t139 10.6405
R8431 DVSS.n312 DVSS.t143 10.6405
R8432 DVSS.n310 DVSS.t142 10.6405
R8433 DVSS.n310 DVSS.t141 10.6405
R8434 DVSS.n112 DVSS.t131 10.6405
R8435 DVSS.n112 DVSS.t127 10.6405
R8436 DVSS.n109 DVSS.t130 10.6405
R8437 DVSS.n109 DVSS.t128 10.6405
R8438 DVSS.n73 DVSS.t89 10.6405
R8439 DVSS.n73 DVSS.t93 10.6405
R8440 DVSS.n72 DVSS.t91 10.6405
R8441 DVSS.n72 DVSS.t92 10.6405
R8442 DVSS.n2579 DVSS.t23 10.6405
R8443 DVSS.n2579 DVSS.t27 10.6405
R8444 DVSS.n2591 DVSS.t26 10.6405
R8445 DVSS.n2591 DVSS.t25 10.6405
R8446 DVSS.n1010 DVSS.n883 10.64
R8447 DVSS.n1192 DVSS.n811 10.64
R8448 DVSS.n1364 DVSS.n610 10.64
R8449 DVSS.n1460 DVSS.n570 10.64
R8450 DVSS.n1536 DVSS.n1535 10.64
R8451 DVSS.n1862 DVSS.n463 10.64
R8452 DVSS.n2044 DVSS.n391 10.64
R8453 DVSS.n2226 DVSS.n319 10.64
R8454 DVSS.n2398 DVSS.n118 10.64
R8455 DVSS.n2494 DVSS.n78 10.64
R8456 DVSS.n2578 DVSS.n2577 10.64
R8457 DVSS.n2768 DVSS.n2761 9.3005
R8458 DVSS.n2769 DVSS.n2768 9.3005
R8459 DVSS.n2735 DVSS.n2734 9.3005
R8460 DVSS.n2735 DVSS.n20 9.3005
R8461 DVSS.n2722 DVSS.n19 9.3005
R8462 DVSS.n2724 DVSS.n19 9.3005
R8463 DVSS.n2741 DVSS.n2740 9.3005
R8464 DVSS.n2740 DVSS.n2739 9.3005
R8465 DVSS.n2684 DVSS.n2680 9.3005
R8466 DVSS.n2685 DVSS.n2684 9.3005
R8467 DVSS.n225 DVSS.n224 9.3005
R8468 DVSS.n224 DVSS.n223 9.3005
R8469 DVSS.n217 DVSS.n216 9.3005
R8470 DVSS.n216 DVSS.n215 9.3005
R8471 DVSS.n2655 DVSS.n2653 9.3005
R8472 DVSS.n2656 DVSS.n2655 9.3005
R8473 DVSS.n248 DVSS.n247 9.3005
R8474 DVSS.n247 DVSS.n244 9.3005
R8475 DVSS.n2359 DVSS.n2358 9.3005
R8476 DVSS.n2359 DVSS.n265 9.3005
R8477 DVSS.n2363 DVSS.n2361 9.3005
R8478 DVSS.n2364 DVSS.n2363 9.3005
R8479 DVSS.n264 DVSS.n140 9.3005
R8480 DVSS.n264 DVSS.n263 9.3005
R8481 DVSS.n2330 DVSS.n2329 9.3005
R8482 DVSS.n2331 DVSS.n2330 9.3005
R8483 DVSS.n2177 DVSS.n2176 9.3005
R8484 DVSS.n2178 DVSS.n2177 9.3005
R8485 DVSS.n2192 DVSS.n2190 9.3005
R8486 DVSS.n2193 DVSS.n2192 9.3005
R8487 DVSS.n2302 DVSS.n2300 9.3005
R8488 DVSS.n2303 DVSS.n2302 9.3005
R8489 DVSS.n2148 DVSS.n2147 9.3005
R8490 DVSS.n2149 DVSS.n2148 9.3005
R8491 DVSS.n1995 DVSS.n1994 9.3005
R8492 DVSS.n1996 DVSS.n1995 9.3005
R8493 DVSS.n2010 DVSS.n2008 9.3005
R8494 DVSS.n2011 DVSS.n2010 9.3005
R8495 DVSS.n2120 DVSS.n2118 9.3005
R8496 DVSS.n2121 DVSS.n2120 9.3005
R8497 DVSS.n1966 DVSS.n1965 9.3005
R8498 DVSS.n1967 DVSS.n1966 9.3005
R8499 DVSS.n1813 DVSS.n1812 9.3005
R8500 DVSS.n1814 DVSS.n1813 9.3005
R8501 DVSS.n1828 DVSS.n1826 9.3005
R8502 DVSS.n1829 DVSS.n1828 9.3005
R8503 DVSS.n1938 DVSS.n1936 9.3005
R8504 DVSS.n1939 DVSS.n1938 9.3005
R8505 DVSS.n1784 DVSS.n1783 9.3005
R8506 DVSS.n1785 DVSS.n1784 9.3005
R8507 DVSS.n1742 DVSS.n1741 9.3005
R8508 DVSS.n1742 DVSS.n512 9.3005
R8509 DVSS.n1729 DVSS.n511 9.3005
R8510 DVSS.n1731 DVSS.n511 9.3005
R8511 DVSS.n1748 DVSS.n1747 9.3005
R8512 DVSS.n1747 DVSS.n1746 9.3005
R8513 DVSS.n1691 DVSS.n1687 9.3005
R8514 DVSS.n1692 DVSS.n1691 9.3005
R8515 DVSS.n717 DVSS.n716 9.3005
R8516 DVSS.n716 DVSS.n715 9.3005
R8517 DVSS.n709 DVSS.n708 9.3005
R8518 DVSS.n708 DVSS.n707 9.3005
R8519 DVSS.n1662 DVSS.n1660 9.3005
R8520 DVSS.n1663 DVSS.n1662 9.3005
R8521 DVSS.n740 DVSS.n739 9.3005
R8522 DVSS.n739 DVSS.n736 9.3005
R8523 DVSS.n1325 DVSS.n1324 9.3005
R8524 DVSS.n1325 DVSS.n757 9.3005
R8525 DVSS.n1329 DVSS.n1327 9.3005
R8526 DVSS.n1330 DVSS.n1329 9.3005
R8527 DVSS.n756 DVSS.n632 9.3005
R8528 DVSS.n756 DVSS.n755 9.3005
R8529 DVSS.n1296 DVSS.n1295 9.3005
R8530 DVSS.n1297 DVSS.n1296 9.3005
R8531 DVSS.n1143 DVSS.n1142 9.3005
R8532 DVSS.n1144 DVSS.n1143 9.3005
R8533 DVSS.n1158 DVSS.n1156 9.3005
R8534 DVSS.n1159 DVSS.n1158 9.3005
R8535 DVSS.n1268 DVSS.n1266 9.3005
R8536 DVSS.n1269 DVSS.n1268 9.3005
R8537 DVSS.n1114 DVSS.n1113 9.3005
R8538 DVSS.n1115 DVSS.n1114 9.3005
R8539 DVSS.n961 DVSS.n960 9.3005
R8540 DVSS.n962 DVSS.n961 9.3005
R8541 DVSS.n976 DVSS.n974 9.3005
R8542 DVSS.n977 DVSS.n976 9.3005
R8543 DVSS.n1086 DVSS.n1084 9.3005
R8544 DVSS.n1087 DVSS.n1086 9.3005
R8545 DVSS.n930 DVSS.n929 9.3005
R8546 DVSS.n919 DVSS.n915 9.3005
R8547 DVSS.n924 DVSS.n920 9.3005
R8548 DVSS.n923 DVSS.n922 9.3005
R8549 DVSS.n921 DVSS.n902 9.3005
R8550 DVSS.n958 DVSS.n957 9.3005
R8551 DVSS.n959 DVSS.n900 9.3005
R8552 DVSS.n984 DVSS.n983 9.3005
R8553 DVSS.n982 DVSS.n901 9.3005
R8554 DVSS.n981 DVSS.n980 9.3005
R8555 DVSS.n979 DVSS.n978 9.3005
R8556 DVSS.n973 DVSS.n971 9.3005
R8557 DVSS.n972 DVSS.n855 9.3005
R8558 DVSS.n1083 DVSS.n1082 9.3005
R8559 DVSS.n1088 DVSS.n853 9.3005
R8560 DVSS.n1091 DVSS.n1090 9.3005
R8561 DVSS.n1089 DVSS.n849 9.3005
R8562 DVSS.n1098 DVSS.n1097 9.3005
R8563 DVSS.n1099 DVSS.n848 9.3005
R8564 DVSS.n1102 DVSS.n1101 9.3005
R8565 DVSS.n1100 DVSS.n843 9.3005
R8566 DVSS.n1111 DVSS.n1110 9.3005
R8567 DVSS.n1112 DVSS.n839 9.3005
R8568 DVSS.n1117 DVSS.n1116 9.3005
R8569 DVSS.n1119 DVSS.n1118 9.3005
R8570 DVSS.n1122 DVSS.n1121 9.3005
R8571 DVSS.n1120 DVSS.n835 9.3005
R8572 DVSS.n1129 DVSS.n1128 9.3005
R8573 DVSS.n1130 DVSS.n834 9.3005
R8574 DVSS.n1133 DVSS.n1132 9.3005
R8575 DVSS.n1131 DVSS.n830 9.3005
R8576 DVSS.n1140 DVSS.n1139 9.3005
R8577 DVSS.n1141 DVSS.n828 9.3005
R8578 DVSS.n1166 DVSS.n1165 9.3005
R8579 DVSS.n1164 DVSS.n829 9.3005
R8580 DVSS.n1163 DVSS.n1162 9.3005
R8581 DVSS.n1161 DVSS.n1160 9.3005
R8582 DVSS.n1155 DVSS.n1153 9.3005
R8583 DVSS.n1154 DVSS.n783 9.3005
R8584 DVSS.n1265 DVSS.n1264 9.3005
R8585 DVSS.n1270 DVSS.n781 9.3005
R8586 DVSS.n1273 DVSS.n1272 9.3005
R8587 DVSS.n1271 DVSS.n777 9.3005
R8588 DVSS.n1280 DVSS.n1279 9.3005
R8589 DVSS.n1281 DVSS.n776 9.3005
R8590 DVSS.n1284 DVSS.n1283 9.3005
R8591 DVSS.n1282 DVSS.n771 9.3005
R8592 DVSS.n1293 DVSS.n1292 9.3005
R8593 DVSS.n1294 DVSS.n767 9.3005
R8594 DVSS.n1299 DVSS.n1298 9.3005
R8595 DVSS.n1301 DVSS.n1300 9.3005
R8596 DVSS.n1304 DVSS.n1303 9.3005
R8597 DVSS.n1302 DVSS.n763 9.3005
R8598 DVSS.n1311 DVSS.n1310 9.3005
R8599 DVSS.n1312 DVSS.n762 9.3005
R8600 DVSS.n1315 DVSS.n1314 9.3005
R8601 DVSS.n1313 DVSS.n758 9.3005
R8602 DVSS.n1322 DVSS.n1321 9.3005
R8603 DVSS.n1323 DVSS.n627 9.3005
R8604 DVSS.n1337 DVSS.n1336 9.3005
R8605 DVSS.n1335 DVSS.n628 9.3005
R8606 DVSS.n1334 DVSS.n1333 9.3005
R8607 DVSS.n1332 DVSS.n1331 9.3005
R8608 DVSS.n660 DVSS.n631 9.3005
R8609 DVSS.n662 DVSS.n661 9.3005
R8610 DVSS.n635 DVSS.n634 9.3005
R8611 DVSS.n754 DVSS.n753 9.3005
R8612 DVSS.n752 DVSS.n751 9.3005
R8613 DVSS.n750 DVSS.n638 9.3005
R8614 DVSS.n749 DVSS.n748 9.3005
R8615 DVSS.n747 DVSS.n746 9.3005
R8616 DVSS.n745 DVSS.n641 9.3005
R8617 DVSS.n744 DVSS.n743 9.3005
R8618 DVSS.n742 DVSS.n741 9.3005
R8619 DVSS.n645 DVSS.n644 9.3005
R8620 DVSS.n735 DVSS.n734 9.3005
R8621 DVSS.n733 DVSS.n732 9.3005
R8622 DVSS.n731 DVSS.n730 9.3005
R8623 DVSS.n729 DVSS.n728 9.3005
R8624 DVSS.n727 DVSS.n650 9.3005
R8625 DVSS.n726 DVSS.n725 9.3005
R8626 DVSS.n724 DVSS.n723 9.3005
R8627 DVSS.n722 DVSS.n653 9.3005
R8628 DVSS.n721 DVSS.n720 9.3005
R8629 DVSS.n719 DVSS.n718 9.3005
R8630 DVSS.n714 DVSS.n656 9.3005
R8631 DVSS.n713 DVSS.n712 9.3005
R8632 DVSS.n711 DVSS.n710 9.3005
R8633 DVSS.n705 DVSS.n703 9.3005
R8634 DVSS.n706 DVSS.n541 9.3005
R8635 DVSS.n1658 DVSS.n1657 9.3005
R8636 DVSS.n1659 DVSS.n539 9.3005
R8637 DVSS.n1666 DVSS.n1665 9.3005
R8638 DVSS.n1664 DVSS.n536 9.3005
R8639 DVSS.n1673 DVSS.n1672 9.3005
R8640 DVSS.n1674 DVSS.n535 9.3005
R8641 DVSS.n1677 DVSS.n1676 9.3005
R8642 DVSS.n1675 DVSS.n531 9.3005
R8643 DVSS.n1685 DVSS.n1684 9.3005
R8644 DVSS.n1686 DVSS.n530 9.3005
R8645 DVSS.n1694 DVSS.n1693 9.3005
R8646 DVSS.n1688 DVSS.n527 9.3005
R8647 DVSS.n1701 DVSS.n1700 9.3005
R8648 DVSS.n1702 DVSS.n526 9.3005
R8649 DVSS.n1705 DVSS.n1704 9.3005
R8650 DVSS.n1703 DVSS.n522 9.3005
R8651 DVSS.n1713 DVSS.n1712 9.3005
R8652 DVSS.n1714 DVSS.n521 9.3005
R8653 DVSS.n1717 DVSS.n1716 9.3005
R8654 DVSS.n1715 DVSS.n513 9.3005
R8655 DVSS.n1740 DVSS.n1739 9.3005
R8656 DVSS.n1738 DVSS.n1737 9.3005
R8657 DVSS.n1736 DVSS.n516 9.3005
R8658 DVSS.n1735 DVSS.n1734 9.3005
R8659 DVSS.n1733 DVSS.n1732 9.3005
R8660 DVSS.n1730 DVSS.n509 9.3005
R8661 DVSS.n1750 DVSS.n1749 9.3005
R8662 DVSS.n1745 DVSS.n505 9.3005
R8663 DVSS.n1758 DVSS.n1757 9.3005
R8664 DVSS.n1759 DVSS.n504 9.3005
R8665 DVSS.n1762 DVSS.n1761 9.3005
R8666 DVSS.n1760 DVSS.n500 9.3005
R8667 DVSS.n1769 DVSS.n1768 9.3005
R8668 DVSS.n1770 DVSS.n499 9.3005
R8669 DVSS.n1773 DVSS.n1772 9.3005
R8670 DVSS.n1771 DVSS.n495 9.3005
R8671 DVSS.n1782 DVSS.n1781 9.3005
R8672 DVSS.n1787 DVSS.n1786 9.3005
R8673 DVSS.n1789 DVSS.n1788 9.3005
R8674 DVSS.n1792 DVSS.n1791 9.3005
R8675 DVSS.n1790 DVSS.n487 9.3005
R8676 DVSS.n1799 DVSS.n1798 9.3005
R8677 DVSS.n1800 DVSS.n486 9.3005
R8678 DVSS.n1803 DVSS.n1802 9.3005
R8679 DVSS.n1801 DVSS.n482 9.3005
R8680 DVSS.n1810 DVSS.n1809 9.3005
R8681 DVSS.n1811 DVSS.n480 9.3005
R8682 DVSS.n1836 DVSS.n1835 9.3005
R8683 DVSS.n1834 DVSS.n481 9.3005
R8684 DVSS.n1833 DVSS.n1832 9.3005
R8685 DVSS.n1831 DVSS.n1830 9.3005
R8686 DVSS.n1825 DVSS.n1823 9.3005
R8687 DVSS.n1824 DVSS.n435 9.3005
R8688 DVSS.n1935 DVSS.n1934 9.3005
R8689 DVSS.n1940 DVSS.n433 9.3005
R8690 DVSS.n1943 DVSS.n1942 9.3005
R8691 DVSS.n1941 DVSS.n429 9.3005
R8692 DVSS.n1950 DVSS.n1949 9.3005
R8693 DVSS.n1951 DVSS.n428 9.3005
R8694 DVSS.n1954 DVSS.n1953 9.3005
R8695 DVSS.n1952 DVSS.n423 9.3005
R8696 DVSS.n1963 DVSS.n1962 9.3005
R8697 DVSS.n1964 DVSS.n419 9.3005
R8698 DVSS.n1969 DVSS.n1968 9.3005
R8699 DVSS.n1971 DVSS.n1970 9.3005
R8700 DVSS.n1974 DVSS.n1973 9.3005
R8701 DVSS.n1972 DVSS.n415 9.3005
R8702 DVSS.n1981 DVSS.n1980 9.3005
R8703 DVSS.n1982 DVSS.n414 9.3005
R8704 DVSS.n1985 DVSS.n1984 9.3005
R8705 DVSS.n1983 DVSS.n410 9.3005
R8706 DVSS.n1992 DVSS.n1991 9.3005
R8707 DVSS.n1993 DVSS.n408 9.3005
R8708 DVSS.n2018 DVSS.n2017 9.3005
R8709 DVSS.n2016 DVSS.n409 9.3005
R8710 DVSS.n2015 DVSS.n2014 9.3005
R8711 DVSS.n2013 DVSS.n2012 9.3005
R8712 DVSS.n2007 DVSS.n2005 9.3005
R8713 DVSS.n2006 DVSS.n363 9.3005
R8714 DVSS.n2117 DVSS.n2116 9.3005
R8715 DVSS.n2122 DVSS.n361 9.3005
R8716 DVSS.n2125 DVSS.n2124 9.3005
R8717 DVSS.n2123 DVSS.n357 9.3005
R8718 DVSS.n2132 DVSS.n2131 9.3005
R8719 DVSS.n2133 DVSS.n356 9.3005
R8720 DVSS.n2136 DVSS.n2135 9.3005
R8721 DVSS.n2134 DVSS.n351 9.3005
R8722 DVSS.n2145 DVSS.n2144 9.3005
R8723 DVSS.n2146 DVSS.n347 9.3005
R8724 DVSS.n2151 DVSS.n2150 9.3005
R8725 DVSS.n2153 DVSS.n2152 9.3005
R8726 DVSS.n2156 DVSS.n2155 9.3005
R8727 DVSS.n2154 DVSS.n343 9.3005
R8728 DVSS.n2163 DVSS.n2162 9.3005
R8729 DVSS.n2164 DVSS.n342 9.3005
R8730 DVSS.n2167 DVSS.n2166 9.3005
R8731 DVSS.n2165 DVSS.n338 9.3005
R8732 DVSS.n2174 DVSS.n2173 9.3005
R8733 DVSS.n2175 DVSS.n336 9.3005
R8734 DVSS.n2200 DVSS.n2199 9.3005
R8735 DVSS.n2198 DVSS.n337 9.3005
R8736 DVSS.n2197 DVSS.n2196 9.3005
R8737 DVSS.n2195 DVSS.n2194 9.3005
R8738 DVSS.n2189 DVSS.n2187 9.3005
R8739 DVSS.n2188 DVSS.n291 9.3005
R8740 DVSS.n2299 DVSS.n2298 9.3005
R8741 DVSS.n2304 DVSS.n289 9.3005
R8742 DVSS.n2307 DVSS.n2306 9.3005
R8743 DVSS.n2305 DVSS.n285 9.3005
R8744 DVSS.n2314 DVSS.n2313 9.3005
R8745 DVSS.n2315 DVSS.n284 9.3005
R8746 DVSS.n2318 DVSS.n2317 9.3005
R8747 DVSS.n2316 DVSS.n279 9.3005
R8748 DVSS.n2327 DVSS.n2326 9.3005
R8749 DVSS.n2328 DVSS.n275 9.3005
R8750 DVSS.n2333 DVSS.n2332 9.3005
R8751 DVSS.n2335 DVSS.n2334 9.3005
R8752 DVSS.n2338 DVSS.n2337 9.3005
R8753 DVSS.n2336 DVSS.n271 9.3005
R8754 DVSS.n2345 DVSS.n2344 9.3005
R8755 DVSS.n2346 DVSS.n270 9.3005
R8756 DVSS.n2349 DVSS.n2348 9.3005
R8757 DVSS.n2347 DVSS.n266 9.3005
R8758 DVSS.n2356 DVSS.n2355 9.3005
R8759 DVSS.n2357 DVSS.n135 9.3005
R8760 DVSS.n2371 DVSS.n2370 9.3005
R8761 DVSS.n2369 DVSS.n136 9.3005
R8762 DVSS.n2368 DVSS.n2367 9.3005
R8763 DVSS.n2366 DVSS.n2365 9.3005
R8764 DVSS.n168 DVSS.n139 9.3005
R8765 DVSS.n170 DVSS.n169 9.3005
R8766 DVSS.n143 DVSS.n142 9.3005
R8767 DVSS.n262 DVSS.n261 9.3005
R8768 DVSS.n260 DVSS.n259 9.3005
R8769 DVSS.n258 DVSS.n146 9.3005
R8770 DVSS.n257 DVSS.n256 9.3005
R8771 DVSS.n255 DVSS.n254 9.3005
R8772 DVSS.n253 DVSS.n149 9.3005
R8773 DVSS.n252 DVSS.n251 9.3005
R8774 DVSS.n250 DVSS.n249 9.3005
R8775 DVSS.n153 DVSS.n152 9.3005
R8776 DVSS.n243 DVSS.n242 9.3005
R8777 DVSS.n241 DVSS.n240 9.3005
R8778 DVSS.n239 DVSS.n238 9.3005
R8779 DVSS.n237 DVSS.n236 9.3005
R8780 DVSS.n235 DVSS.n158 9.3005
R8781 DVSS.n234 DVSS.n233 9.3005
R8782 DVSS.n232 DVSS.n231 9.3005
R8783 DVSS.n230 DVSS.n161 9.3005
R8784 DVSS.n229 DVSS.n228 9.3005
R8785 DVSS.n227 DVSS.n226 9.3005
R8786 DVSS.n222 DVSS.n164 9.3005
R8787 DVSS.n221 DVSS.n220 9.3005
R8788 DVSS.n219 DVSS.n218 9.3005
R8789 DVSS.n213 DVSS.n211 9.3005
R8790 DVSS.n214 DVSS.n49 9.3005
R8791 DVSS.n2651 DVSS.n2650 9.3005
R8792 DVSS.n2652 DVSS.n47 9.3005
R8793 DVSS.n2659 DVSS.n2658 9.3005
R8794 DVSS.n2657 DVSS.n44 9.3005
R8795 DVSS.n2666 DVSS.n2665 9.3005
R8796 DVSS.n2667 DVSS.n43 9.3005
R8797 DVSS.n2670 DVSS.n2669 9.3005
R8798 DVSS.n2668 DVSS.n39 9.3005
R8799 DVSS.n2678 DVSS.n2677 9.3005
R8800 DVSS.n2679 DVSS.n38 9.3005
R8801 DVSS.n2687 DVSS.n2686 9.3005
R8802 DVSS.n2681 DVSS.n35 9.3005
R8803 DVSS.n2694 DVSS.n2693 9.3005
R8804 DVSS.n2695 DVSS.n34 9.3005
R8805 DVSS.n2698 DVSS.n2697 9.3005
R8806 DVSS.n2696 DVSS.n30 9.3005
R8807 DVSS.n2706 DVSS.n2705 9.3005
R8808 DVSS.n2707 DVSS.n29 9.3005
R8809 DVSS.n2710 DVSS.n2709 9.3005
R8810 DVSS.n2708 DVSS.n21 9.3005
R8811 DVSS.n2733 DVSS.n2732 9.3005
R8812 DVSS.n2731 DVSS.n2730 9.3005
R8813 DVSS.n2729 DVSS.n24 9.3005
R8814 DVSS.n2728 DVSS.n2727 9.3005
R8815 DVSS.n2726 DVSS.n2725 9.3005
R8816 DVSS.n2723 DVSS.n17 9.3005
R8817 DVSS.n2743 DVSS.n2742 9.3005
R8818 DVSS.n2738 DVSS.n13 9.3005
R8819 DVSS.n2751 DVSS.n2750 9.3005
R8820 DVSS.n2752 DVSS.n11 9.3005
R8821 DVSS.n2781 DVSS.n2780 9.3005
R8822 DVSS.n2779 DVSS.n12 9.3005
R8823 DVSS.n2778 DVSS.n2777 9.3005
R8824 DVSS.n2776 DVSS.n2775 9.3005
R8825 DVSS.n2774 DVSS.n2755 9.3005
R8826 DVSS.n2773 DVSS.n2772 9.3005
R8827 DVSS.n2771 DVSS.n2770 9.3005
R8828 DVSS.n2765 DVSS.n2760 9.3005
R8829 DVSS.n2764 DVSS.n2763 9.3005
R8830 DVSS.n2620 DVSS.n2619 9.3005
R8831 DVSS.n2617 DVSS.n2616 9.3005
R8832 DVSS.n2593 DVSS.n2592 9.3005
R8833 DVSS.n2610 DVSS.n2609 9.3005
R8834 DVSS.n2609 DVSS.n2608 9.3005
R8835 DVSS.n2631 DVSS.n2630 9.3005
R8836 DVSS.n2571 DVSS.n2560 9.3005
R8837 DVSS.n2543 DVSS.n2542 9.3005
R8838 DVSS.n2544 DVSS.n63 9.3005
R8839 DVSS.n2546 DVSS.n2545 9.3005
R8840 DVSS.n2497 DVSS.n2496 9.3005
R8841 DVSS.n2500 DVSS.n2499 9.3005
R8842 DVSS.n2513 DVSS.n2512 9.3005
R8843 DVSS.n2518 DVSS.n2517 9.3005
R8844 DVSS.n2517 DVSS.n2516 9.3005
R8845 DVSS.n2480 DVSS.n83 9.3005
R8846 DVSS.n2484 DVSS.n2483 9.3005
R8847 DVSS.n2449 DVSS.n99 9.3005
R8848 DVSS.n2451 DVSS.n2450 9.3005
R8849 DVSS.n2453 DVSS.n2452 9.3005
R8850 DVSS.n2411 DVSS.n2410 9.3005
R8851 DVSS.n2414 DVSS.n2413 9.3005
R8852 DVSS.n2428 DVSS.n2427 9.3005
R8853 DVSS.n2430 DVSS.n111 9.3005
R8854 DVSS.n2431 DVSS.n2430 9.3005
R8855 DVSS.n2392 DVSS.n123 9.3005
R8856 DVSS.n2396 DVSS.n2395 9.3005
R8857 DVSS.n2277 DVSS.n2276 9.3005
R8858 DVSS.n2280 DVSS.n2279 9.3005
R8859 DVSS.n2278 DVSS.n300 9.3005
R8860 DVSS.n2239 DVSS.n2238 9.3005
R8861 DVSS.n2242 DVSS.n2241 9.3005
R8862 DVSS.n2253 DVSS.n2252 9.3005
R8863 DVSS.n2255 DVSS.n311 9.3005
R8864 DVSS.n2256 DVSS.n2255 9.3005
R8865 DVSS.n2220 DVSS.n324 9.3005
R8866 DVSS.n2224 DVSS.n2223 9.3005
R8867 DVSS.n2095 DVSS.n2094 9.3005
R8868 DVSS.n2098 DVSS.n2097 9.3005
R8869 DVSS.n2096 DVSS.n372 9.3005
R8870 DVSS.n2057 DVSS.n2056 9.3005
R8871 DVSS.n2060 DVSS.n2059 9.3005
R8872 DVSS.n2071 DVSS.n2070 9.3005
R8873 DVSS.n2073 DVSS.n383 9.3005
R8874 DVSS.n2074 DVSS.n2073 9.3005
R8875 DVSS.n2038 DVSS.n396 9.3005
R8876 DVSS.n2042 DVSS.n2041 9.3005
R8877 DVSS.n1913 DVSS.n1912 9.3005
R8878 DVSS.n1916 DVSS.n1915 9.3005
R8879 DVSS.n1914 DVSS.n444 9.3005
R8880 DVSS.n1875 DVSS.n1874 9.3005
R8881 DVSS.n1878 DVSS.n1877 9.3005
R8882 DVSS.n1889 DVSS.n1888 9.3005
R8883 DVSS.n1891 DVSS.n455 9.3005
R8884 DVSS.n1892 DVSS.n1891 9.3005
R8885 DVSS.n1856 DVSS.n468 9.3005
R8886 DVSS.n1860 DVSS.n1859 9.3005
R8887 DVSS.n1602 DVSS.n1601 9.3005
R8888 DVSS.n1600 DVSS.n1558 9.3005
R8889 DVSS.n1560 DVSS.n1559 9.3005
R8890 DVSS.n1627 DVSS.n1626 9.3005
R8891 DVSS.n1624 DVSS.n1623 9.3005
R8892 DVSS.n1547 DVSS.n1546 9.3005
R8893 DVSS.n1617 DVSS.n1616 9.3005
R8894 DVSS.n1616 DVSS.n1615 9.3005
R8895 DVSS.n1638 DVSS.n1637 9.3005
R8896 DVSS.n1531 DVSS.n1526 9.3005
R8897 DVSS.n1509 DVSS.n1508 9.3005
R8898 DVSS.n1510 DVSS.n555 9.3005
R8899 DVSS.n1512 DVSS.n1511 9.3005
R8900 DVSS.n1463 DVSS.n1462 9.3005
R8901 DVSS.n1466 DVSS.n1465 9.3005
R8902 DVSS.n1479 DVSS.n1478 9.3005
R8903 DVSS.n1484 DVSS.n1483 9.3005
R8904 DVSS.n1483 DVSS.n1482 9.3005
R8905 DVSS.n1446 DVSS.n575 9.3005
R8906 DVSS.n1450 DVSS.n1449 9.3005
R8907 DVSS.n1415 DVSS.n591 9.3005
R8908 DVSS.n1417 DVSS.n1416 9.3005
R8909 DVSS.n1419 DVSS.n1418 9.3005
R8910 DVSS.n1377 DVSS.n1376 9.3005
R8911 DVSS.n1380 DVSS.n1379 9.3005
R8912 DVSS.n1394 DVSS.n1393 9.3005
R8913 DVSS.n1396 DVSS.n603 9.3005
R8914 DVSS.n1397 DVSS.n1396 9.3005
R8915 DVSS.n1358 DVSS.n615 9.3005
R8916 DVSS.n1362 DVSS.n1361 9.3005
R8917 DVSS.n1243 DVSS.n1242 9.3005
R8918 DVSS.n1246 DVSS.n1245 9.3005
R8919 DVSS.n1244 DVSS.n792 9.3005
R8920 DVSS.n1205 DVSS.n1204 9.3005
R8921 DVSS.n1208 DVSS.n1207 9.3005
R8922 DVSS.n1219 DVSS.n1218 9.3005
R8923 DVSS.n1221 DVSS.n803 9.3005
R8924 DVSS.n1222 DVSS.n1221 9.3005
R8925 DVSS.n1186 DVSS.n816 9.3005
R8926 DVSS.n1190 DVSS.n1189 9.3005
R8927 DVSS.n1061 DVSS.n1060 9.3005
R8928 DVSS.n1064 DVSS.n1063 9.3005
R8929 DVSS.n1062 DVSS.n864 9.3005
R8930 DVSS.n1023 DVSS.n1022 9.3005
R8931 DVSS.n1026 DVSS.n1025 9.3005
R8932 DVSS.n1037 DVSS.n1036 9.3005
R8933 DVSS.n1039 DVSS.n875 9.3005
R8934 DVSS.n1040 DVSS.n1039 9.3005
R8935 DVSS.n1004 DVSS.n888 9.3005
R8936 DVSS.n1008 DVSS.n1007 9.3005
R8937 DVSS.n938 DVSS.n937 9.3005
R8938 DVSS.n941 DVSS.n940 9.3005
R8939 DVSS.n939 DVSS.n909 9.3005
R8940 DVSS.n2787 DVSS.n2786 9.3005
R8941 DVSS.n2603 DVSS.n0 9.3005
R8942 DVSS.n2605 DVSS.n2604 9.3005
R8943 DVSS.n2607 DVSS.n2606 9.3005
R8944 DVSS.n2596 DVSS.n2595 9.3005
R8945 DVSS.n2611 DVSS.n2590 9.3005
R8946 DVSS.n2613 DVSS.n2612 9.3005
R8947 DVSS.n2615 DVSS.n2614 9.3005
R8948 DVSS.n2583 DVSS.n2582 9.3005
R8949 DVSS.n2581 DVSS.n2576 9.3005
R8950 DVSS.n2622 DVSS.n2621 9.3005
R8951 DVSS.n2624 DVSS.n2623 9.3005
R8952 DVSS.n2625 DVSS.n2570 9.3005
R8953 DVSS.n2627 DVSS.n2626 9.3005
R8954 DVSS.n2629 DVSS.n2628 9.3005
R8955 DVSS.n2634 DVSS.n2559 9.3005
R8956 DVSS.n2636 DVSS.n2635 9.3005
R8957 DVSS.n2638 DVSS.n2637 9.3005
R8958 DVSS.n2639 DVSS.n59 9.3005
R8959 DVSS.n2641 DVSS.n2640 9.3005
R8960 DVSS.n2556 DVSS.n58 9.3005
R8961 DVSS.n2555 DVSS.n2554 9.3005
R8962 DVSS.n64 DVSS.n60 9.3005
R8963 DVSS.n2548 DVSS.n2547 9.3005
R8964 DVSS.n2541 DVSS.n62 9.3005
R8965 DVSS.n2538 DVSS.n2537 9.3005
R8966 DVSS.n2529 DVSS.n66 9.3005
R8967 DVSS.n2531 DVSS.n2530 9.3005
R8968 DVSS.n2528 DVSS.n68 9.3005
R8969 DVSS.n2527 DVSS.n2526 9.3005
R8970 DVSS.n2515 DVSS.n69 9.3005
R8971 DVSS.n2520 DVSS.n2519 9.3005
R8972 DVSS.n2511 DVSS.n71 9.3005
R8973 DVSS.n2510 DVSS.n2509 9.3005
R8974 DVSS.n2501 DVSS.n75 9.3005
R8975 DVSS.n2503 DVSS.n2502 9.3005
R8976 DVSS.n2495 DVSS.n77 9.3005
R8977 DVSS.n2493 DVSS.n2492 9.3005
R8978 DVSS.n2485 DVSS.n79 9.3005
R8979 DVSS.n2487 DVSS.n2486 9.3005
R8980 DVSS.n2479 DVSS.n81 9.3005
R8981 DVSS.n2478 DVSS.n2477 9.3005
R8982 DVSS.n2468 DVSS.n84 9.3005
R8983 DVSS.n2470 DVSS.n2469 9.3005
R8984 DVSS.n2467 DVSS.n88 9.3005
R8985 DVSS.n2466 DVSS.n2465 9.3005
R8986 DVSS.n2455 DVSS.n89 9.3005
R8987 DVSS.n2457 DVSS.n2456 9.3005
R8988 DVSS.n2454 DVSS.n97 9.3005
R8989 DVSS.n2446 DVSS.n98 9.3005
R8990 DVSS.n2448 DVSS.n2447 9.3005
R8991 DVSS.n2443 DVSS.n2442 9.3005
R8992 DVSS.n2441 DVSS.n103 9.3005
R8993 DVSS.n2440 DVSS.n2439 9.3005
R8994 DVSS.n2432 DVSS.n106 9.3005
R8995 DVSS.n2434 DVSS.n2433 9.3005
R8996 DVSS.n110 DVSS.n108 9.3005
R8997 DVSS.n2424 DVSS.n2423 9.3005
R8998 DVSS.n2426 DVSS.n2425 9.3005
R8999 DVSS.n117 DVSS.n114 9.3005
R9000 DVSS.n2416 DVSS.n2415 9.3005
R9001 DVSS.n2409 DVSS.n116 9.3005
R9002 DVSS.n2408 DVSS.n2407 9.3005
R9003 DVSS.n2399 DVSS.n119 9.3005
R9004 DVSS.n2401 DVSS.n2400 9.3005
R9005 DVSS.n2397 DVSS.n121 9.3005
R9006 DVSS.n2391 DVSS.n2390 9.3005
R9007 DVSS.n2381 DVSS.n124 9.3005
R9008 DVSS.n2383 DVSS.n2382 9.3005
R9009 DVSS.n2380 DVSS.n128 9.3005
R9010 DVSS.n2379 DVSS.n2378 9.3005
R9011 DVSS.n2287 DVSS.n129 9.3005
R9012 DVSS.n2289 DVSS.n2288 9.3005
R9013 DVSS.n2286 DVSS.n299 9.3005
R9014 DVSS.n2285 DVSS.n2284 9.3005
R9015 DVSS.n2282 DVSS.n2281 9.3005
R9016 DVSS.n2275 DVSS.n301 9.3005
R9017 DVSS.n2272 DVSS.n2271 9.3005
R9018 DVSS.n2268 DVSS.n2267 9.3005
R9019 DVSS.n2266 DVSS.n305 9.3005
R9020 DVSS.n2265 DVSS.n2264 9.3005
R9021 DVSS.n309 DVSS.n306 9.3005
R9022 DVSS.n2258 DVSS.n2257 9.3005
R9023 DVSS.n314 DVSS.n308 9.3005
R9024 DVSS.n2251 DVSS.n2250 9.3005
R9025 DVSS.n318 DVSS.n315 9.3005
R9026 DVSS.n2244 DVSS.n2243 9.3005
R9027 DVSS.n2237 DVSS.n317 9.3005
R9028 DVSS.n2236 DVSS.n2235 9.3005
R9029 DVSS.n2227 DVSS.n320 9.3005
R9030 DVSS.n2229 DVSS.n2228 9.3005
R9031 DVSS.n2225 DVSS.n322 9.3005
R9032 DVSS.n2219 DVSS.n2218 9.3005
R9033 DVSS.n2210 DVSS.n325 9.3005
R9034 DVSS.n2212 DVSS.n2211 9.3005
R9035 DVSS.n2209 DVSS.n329 9.3005
R9036 DVSS.n2208 DVSS.n2207 9.3005
R9037 DVSS.n2105 DVSS.n330 9.3005
R9038 DVSS.n2107 DVSS.n2106 9.3005
R9039 DVSS.n2104 DVSS.n371 9.3005
R9040 DVSS.n2103 DVSS.n2102 9.3005
R9041 DVSS.n2100 DVSS.n2099 9.3005
R9042 DVSS.n2093 DVSS.n373 9.3005
R9043 DVSS.n2090 DVSS.n2089 9.3005
R9044 DVSS.n2086 DVSS.n2085 9.3005
R9045 DVSS.n2084 DVSS.n377 9.3005
R9046 DVSS.n2083 DVSS.n2082 9.3005
R9047 DVSS.n381 DVSS.n378 9.3005
R9048 DVSS.n2076 DVSS.n2075 9.3005
R9049 DVSS.n386 DVSS.n380 9.3005
R9050 DVSS.n2069 DVSS.n2068 9.3005
R9051 DVSS.n390 DVSS.n387 9.3005
R9052 DVSS.n2062 DVSS.n2061 9.3005
R9053 DVSS.n2055 DVSS.n389 9.3005
R9054 DVSS.n2054 DVSS.n2053 9.3005
R9055 DVSS.n2045 DVSS.n392 9.3005
R9056 DVSS.n2047 DVSS.n2046 9.3005
R9057 DVSS.n2043 DVSS.n394 9.3005
R9058 DVSS.n2037 DVSS.n2036 9.3005
R9059 DVSS.n2028 DVSS.n397 9.3005
R9060 DVSS.n2030 DVSS.n2029 9.3005
R9061 DVSS.n2027 DVSS.n401 9.3005
R9062 DVSS.n2026 DVSS.n2025 9.3005
R9063 DVSS.n1923 DVSS.n402 9.3005
R9064 DVSS.n1925 DVSS.n1924 9.3005
R9065 DVSS.n1922 DVSS.n443 9.3005
R9066 DVSS.n1921 DVSS.n1920 9.3005
R9067 DVSS.n1918 DVSS.n1917 9.3005
R9068 DVSS.n1911 DVSS.n445 9.3005
R9069 DVSS.n1908 DVSS.n1907 9.3005
R9070 DVSS.n1904 DVSS.n1903 9.3005
R9071 DVSS.n1902 DVSS.n449 9.3005
R9072 DVSS.n1901 DVSS.n1900 9.3005
R9073 DVSS.n453 DVSS.n450 9.3005
R9074 DVSS.n1894 DVSS.n1893 9.3005
R9075 DVSS.n458 DVSS.n452 9.3005
R9076 DVSS.n1887 DVSS.n1886 9.3005
R9077 DVSS.n462 DVSS.n459 9.3005
R9078 DVSS.n1880 DVSS.n1879 9.3005
R9079 DVSS.n1873 DVSS.n461 9.3005
R9080 DVSS.n1872 DVSS.n1871 9.3005
R9081 DVSS.n1863 DVSS.n464 9.3005
R9082 DVSS.n1865 DVSS.n1864 9.3005
R9083 DVSS.n1861 DVSS.n466 9.3005
R9084 DVSS.n1855 DVSS.n1854 9.3005
R9085 DVSS.n1846 DVSS.n469 9.3005
R9086 DVSS.n1848 DVSS.n1847 9.3005
R9087 DVSS.n1845 DVSS.n473 9.3005
R9088 DVSS.n1844 DVSS.n1843 9.3005
R9089 DVSS.n1564 DVSS.n474 9.3005
R9090 DVSS.n1594 DVSS.n1593 9.3005
R9091 DVSS.n1595 DVSS.n1563 9.3005
R9092 DVSS.n1597 DVSS.n1596 9.3005
R9093 DVSS.n1599 DVSS.n1598 9.3005
R9094 DVSS.n1557 DVSS.n1556 9.3005
R9095 DVSS.n1607 DVSS.n1606 9.3005
R9096 DVSS.n1609 DVSS.n1608 9.3005
R9097 DVSS.n1610 DVSS.n1553 9.3005
R9098 DVSS.n1612 DVSS.n1611 9.3005
R9099 DVSS.n1614 DVSS.n1613 9.3005
R9100 DVSS.n1550 DVSS.n1549 9.3005
R9101 DVSS.n1618 DVSS.n1544 9.3005
R9102 DVSS.n1620 DVSS.n1619 9.3005
R9103 DVSS.n1622 DVSS.n1621 9.3005
R9104 DVSS.n1541 DVSS.n1540 9.3005
R9105 DVSS.n1539 DVSS.n1534 9.3005
R9106 DVSS.n1629 DVSS.n1628 9.3005
R9107 DVSS.n1631 DVSS.n1630 9.3005
R9108 DVSS.n1632 DVSS.n1530 9.3005
R9109 DVSS.n1634 DVSS.n1633 9.3005
R9110 DVSS.n1636 DVSS.n1635 9.3005
R9111 DVSS.n1641 DVSS.n1525 9.3005
R9112 DVSS.n1643 DVSS.n1642 9.3005
R9113 DVSS.n1645 DVSS.n1644 9.3005
R9114 DVSS.n1646 DVSS.n551 9.3005
R9115 DVSS.n1648 DVSS.n1647 9.3005
R9116 DVSS.n1522 DVSS.n550 9.3005
R9117 DVSS.n1521 DVSS.n1520 9.3005
R9118 DVSS.n556 DVSS.n552 9.3005
R9119 DVSS.n1514 DVSS.n1513 9.3005
R9120 DVSS.n1507 DVSS.n554 9.3005
R9121 DVSS.n1504 DVSS.n1503 9.3005
R9122 DVSS.n1495 DVSS.n558 9.3005
R9123 DVSS.n1497 DVSS.n1496 9.3005
R9124 DVSS.n1494 DVSS.n560 9.3005
R9125 DVSS.n1493 DVSS.n1492 9.3005
R9126 DVSS.n1481 DVSS.n561 9.3005
R9127 DVSS.n1486 DVSS.n1485 9.3005
R9128 DVSS.n1477 DVSS.n563 9.3005
R9129 DVSS.n1476 DVSS.n1475 9.3005
R9130 DVSS.n1467 DVSS.n567 9.3005
R9131 DVSS.n1469 DVSS.n1468 9.3005
R9132 DVSS.n1461 DVSS.n569 9.3005
R9133 DVSS.n1459 DVSS.n1458 9.3005
R9134 DVSS.n1451 DVSS.n571 9.3005
R9135 DVSS.n1453 DVSS.n1452 9.3005
R9136 DVSS.n1445 DVSS.n573 9.3005
R9137 DVSS.n1444 DVSS.n1443 9.3005
R9138 DVSS.n1434 DVSS.n576 9.3005
R9139 DVSS.n1436 DVSS.n1435 9.3005
R9140 DVSS.n1433 DVSS.n580 9.3005
R9141 DVSS.n1432 DVSS.n1431 9.3005
R9142 DVSS.n1421 DVSS.n581 9.3005
R9143 DVSS.n1423 DVSS.n1422 9.3005
R9144 DVSS.n1420 DVSS.n589 9.3005
R9145 DVSS.n1412 DVSS.n590 9.3005
R9146 DVSS.n1414 DVSS.n1413 9.3005
R9147 DVSS.n1409 DVSS.n1408 9.3005
R9148 DVSS.n1407 DVSS.n595 9.3005
R9149 DVSS.n1406 DVSS.n1405 9.3005
R9150 DVSS.n1398 DVSS.n598 9.3005
R9151 DVSS.n1400 DVSS.n1399 9.3005
R9152 DVSS.n602 DVSS.n600 9.3005
R9153 DVSS.n1390 DVSS.n1389 9.3005
R9154 DVSS.n1392 DVSS.n1391 9.3005
R9155 DVSS.n609 DVSS.n606 9.3005
R9156 DVSS.n1382 DVSS.n1381 9.3005
R9157 DVSS.n1375 DVSS.n608 9.3005
R9158 DVSS.n1374 DVSS.n1373 9.3005
R9159 DVSS.n1365 DVSS.n611 9.3005
R9160 DVSS.n1367 DVSS.n1366 9.3005
R9161 DVSS.n1363 DVSS.n613 9.3005
R9162 DVSS.n1357 DVSS.n1356 9.3005
R9163 DVSS.n1347 DVSS.n616 9.3005
R9164 DVSS.n1349 DVSS.n1348 9.3005
R9165 DVSS.n1346 DVSS.n620 9.3005
R9166 DVSS.n1345 DVSS.n1344 9.3005
R9167 DVSS.n1253 DVSS.n621 9.3005
R9168 DVSS.n1255 DVSS.n1254 9.3005
R9169 DVSS.n1252 DVSS.n791 9.3005
R9170 DVSS.n1251 DVSS.n1250 9.3005
R9171 DVSS.n1248 DVSS.n1247 9.3005
R9172 DVSS.n1241 DVSS.n793 9.3005
R9173 DVSS.n1238 DVSS.n1237 9.3005
R9174 DVSS.n1234 DVSS.n1233 9.3005
R9175 DVSS.n1232 DVSS.n797 9.3005
R9176 DVSS.n1231 DVSS.n1230 9.3005
R9177 DVSS.n801 DVSS.n798 9.3005
R9178 DVSS.n1224 DVSS.n1223 9.3005
R9179 DVSS.n806 DVSS.n800 9.3005
R9180 DVSS.n1217 DVSS.n1216 9.3005
R9181 DVSS.n810 DVSS.n807 9.3005
R9182 DVSS.n1210 DVSS.n1209 9.3005
R9183 DVSS.n1203 DVSS.n809 9.3005
R9184 DVSS.n1202 DVSS.n1201 9.3005
R9185 DVSS.n1193 DVSS.n812 9.3005
R9186 DVSS.n1195 DVSS.n1194 9.3005
R9187 DVSS.n1191 DVSS.n814 9.3005
R9188 DVSS.n1185 DVSS.n1184 9.3005
R9189 DVSS.n1176 DVSS.n817 9.3005
R9190 DVSS.n1178 DVSS.n1177 9.3005
R9191 DVSS.n1175 DVSS.n821 9.3005
R9192 DVSS.n1174 DVSS.n1173 9.3005
R9193 DVSS.n1071 DVSS.n822 9.3005
R9194 DVSS.n1073 DVSS.n1072 9.3005
R9195 DVSS.n1070 DVSS.n863 9.3005
R9196 DVSS.n1069 DVSS.n1068 9.3005
R9197 DVSS.n1066 DVSS.n1065 9.3005
R9198 DVSS.n1059 DVSS.n865 9.3005
R9199 DVSS.n1056 DVSS.n1055 9.3005
R9200 DVSS.n1052 DVSS.n1051 9.3005
R9201 DVSS.n1050 DVSS.n869 9.3005
R9202 DVSS.n1049 DVSS.n1048 9.3005
R9203 DVSS.n873 DVSS.n870 9.3005
R9204 DVSS.n1042 DVSS.n1041 9.3005
R9205 DVSS.n878 DVSS.n872 9.3005
R9206 DVSS.n1035 DVSS.n1034 9.3005
R9207 DVSS.n882 DVSS.n879 9.3005
R9208 DVSS.n1028 DVSS.n1027 9.3005
R9209 DVSS.n1021 DVSS.n881 9.3005
R9210 DVSS.n1020 DVSS.n1019 9.3005
R9211 DVSS.n1011 DVSS.n884 9.3005
R9212 DVSS.n1013 DVSS.n1012 9.3005
R9213 DVSS.n1009 DVSS.n886 9.3005
R9214 DVSS.n1003 DVSS.n1002 9.3005
R9215 DVSS.n994 DVSS.n889 9.3005
R9216 DVSS.n996 DVSS.n995 9.3005
R9217 DVSS.n993 DVSS.n893 9.3005
R9218 DVSS.n992 DVSS.n991 9.3005
R9219 DVSS.n948 DVSS.n894 9.3005
R9220 DVSS.n950 DVSS.n949 9.3005
R9221 DVSS.n947 DVSS.n908 9.3005
R9222 DVSS.n946 DVSS.n945 9.3005
R9223 DVSS.n943 DVSS.n942 9.3005
R9224 DVSS.n936 DVSS.n910 9.3005
R9225 DVSS.n933 DVSS.n932 9.3005
R9226 DVSS.n1114 DVSS.n842 8.54791
R9227 DVSS.n1296 DVSS.n770 8.54791
R9228 DVSS.n739 DVSS.n738 8.54791
R9229 DVSS.n1691 DVSS.n1690 8.54791
R9230 DVSS.n1784 DVSS.n494 8.54791
R9231 DVSS.n1966 DVSS.n422 8.54791
R9232 DVSS.n2148 DVSS.n350 8.54791
R9233 DVSS.n2330 DVSS.n278 8.54791
R9234 DVSS.n247 DVSS.n246 8.54791
R9235 DVSS.n2684 DVSS.n2683 8.54791
R9236 DVSS.n2768 DVSS.n2767 8.54791
R9237 DVSS.n842 DVSS 8.43944
R9238 DVSS.n770 DVSS 8.43944
R9239 DVSS.n738 DVSS 8.43944
R9240 DVSS.n1690 DVSS 8.43944
R9241 DVSS.n494 DVSS 8.43944
R9242 DVSS.n422 DVSS 8.43944
R9243 DVSS.n350 DVSS 8.43944
R9244 DVSS.n278 DVSS 8.43944
R9245 DVSS.n246 DVSS 8.43944
R9246 DVSS.n2683 DVSS 8.43944
R9247 DVSS.n2767 DVSS 8.43944
R9248 DVSS.n1007 DVSS 6.4005
R9249 DVSS.n1189 DVSS 6.4005
R9250 DVSS.n1361 DVSS 6.4005
R9251 DVSS.n1449 DVSS 6.4005
R9252 DVSS.n1526 DVSS 6.4005
R9253 DVSS.n1859 DVSS 6.4005
R9254 DVSS.n2041 DVSS 6.4005
R9255 DVSS.n2223 DVSS 6.4005
R9256 DVSS.n2395 DVSS 6.4005
R9257 DVSS.n2483 DVSS 6.4005
R9258 DVSS.n2560 DVSS 6.4005
R9259 DVSS.n940 DVSS.n938 6.36434
R9260 DVSS.n1063 DVSS.n1061 6.36434
R9261 DVSS.n1245 DVSS.n1243 6.36434
R9262 DVSS.n1417 DVSS.n591 6.36434
R9263 DVSS.n1510 DVSS.n1509 6.36434
R9264 DVSS.n1602 DVSS.n1558 6.36434
R9265 DVSS.n1915 DVSS.n1913 6.36434
R9266 DVSS.n2097 DVSS.n2095 6.36434
R9267 DVSS.n2279 DVSS.n2277 6.36434
R9268 DVSS.n2451 DVSS.n99 6.36434
R9269 DVSS.n2544 DVSS.n2543 6.36434
R9270 DVSS.n940 DVSS.n939 6.00276
R9271 DVSS.n1063 DVSS.n1062 6.00276
R9272 DVSS.n1245 DVSS.n1244 6.00276
R9273 DVSS.n1418 DVSS.n1417 6.00276
R9274 DVSS.n1511 DVSS.n1510 6.00276
R9275 DVSS.n1559 DVSS.n1558 6.00276
R9276 DVSS.n1915 DVSS.n1914 6.00276
R9277 DVSS.n2097 DVSS.n2096 6.00276
R9278 DVSS.n2279 DVSS.n2278 6.00276
R9279 DVSS.n2452 DVSS.n2451 6.00276
R9280 DVSS.n2545 DVSS.n2544 6.00276
R9281 DVSS.n931 DVSS.n914 5.46185
R9282 DVSS.n1006 DVSS 5.45235
R9283 DVSS.n1188 DVSS 5.45235
R9284 DVSS.n1360 DVSS 5.45235
R9285 DVSS.n1448 DVSS 5.45235
R9286 DVSS.n1639 DVSS 5.45235
R9287 DVSS.n1858 DVSS 5.45235
R9288 DVSS.n2040 DVSS 5.45235
R9289 DVSS.n2222 DVSS 5.45235
R9290 DVSS.n2394 DVSS 5.45235
R9291 DVSS.n2482 DVSS 5.45235
R9292 DVSS.n2632 DVSS 5.45235
R9293 DVSS.n929 DVSS.n914 4.06937
R9294 DVSS.n929 DVSS.n915 4.06937
R9295 DVSS.n924 DVSS.n915 4.06937
R9296 DVSS.n924 DVSS.n923 4.06937
R9297 DVSS.n923 DVSS.n902 4.06937
R9298 DVSS.n957 DVSS.n902 4.06937
R9299 DVSS.n957 DVSS.n900 4.06937
R9300 DVSS.n984 DVSS.n900 4.06937
R9301 DVSS.n984 DVSS.n901 4.06937
R9302 DVSS.n980 DVSS.n901 4.06937
R9303 DVSS.n980 DVSS.n979 4.06937
R9304 DVSS.n979 DVSS.n971 4.06937
R9305 DVSS.n971 DVSS.n855 4.06937
R9306 DVSS.n1082 DVSS.n855 4.06937
R9307 DVSS.n1082 DVSS.n853 4.06937
R9308 DVSS.n1091 DVSS.n853 4.06937
R9309 DVSS.n1091 DVSS.n849 4.06937
R9310 DVSS.n1097 DVSS.n849 4.06937
R9311 DVSS.n1097 DVSS.n848 4.06937
R9312 DVSS.n1102 DVSS.n848 4.06937
R9313 DVSS.n1102 DVSS.n843 4.06937
R9314 DVSS.n1110 DVSS.n843 4.06937
R9315 DVSS.n1110 DVSS.n839 4.06937
R9316 DVSS.n1117 DVSS.n839 4.06937
R9317 DVSS.n1118 DVSS.n1117 4.06937
R9318 DVSS.n1122 DVSS.n835 4.06937
R9319 DVSS.n1128 DVSS.n835 4.06937
R9320 DVSS.n1128 DVSS.n834 4.06937
R9321 DVSS.n1133 DVSS.n834 4.06937
R9322 DVSS.n1133 DVSS.n830 4.06937
R9323 DVSS.n1139 DVSS.n830 4.06937
R9324 DVSS.n1139 DVSS.n828 4.06937
R9325 DVSS.n1166 DVSS.n828 4.06937
R9326 DVSS.n1166 DVSS.n829 4.06937
R9327 DVSS.n1162 DVSS.n829 4.06937
R9328 DVSS.n1162 DVSS.n1161 4.06937
R9329 DVSS.n1161 DVSS.n1153 4.06937
R9330 DVSS.n1153 DVSS.n783 4.06937
R9331 DVSS.n1264 DVSS.n783 4.06937
R9332 DVSS.n1264 DVSS.n781 4.06937
R9333 DVSS.n1273 DVSS.n781 4.06937
R9334 DVSS.n1273 DVSS.n777 4.06937
R9335 DVSS.n1279 DVSS.n777 4.06937
R9336 DVSS.n1279 DVSS.n776 4.06937
R9337 DVSS.n1284 DVSS.n776 4.06937
R9338 DVSS.n1284 DVSS.n771 4.06937
R9339 DVSS.n1292 DVSS.n771 4.06937
R9340 DVSS.n1292 DVSS.n767 4.06937
R9341 DVSS.n1299 DVSS.n767 4.06937
R9342 DVSS.n1300 DVSS.n1299 4.06937
R9343 DVSS.n1304 DVSS.n763 4.06937
R9344 DVSS.n1310 DVSS.n763 4.06937
R9345 DVSS.n1310 DVSS.n762 4.06937
R9346 DVSS.n1315 DVSS.n762 4.06937
R9347 DVSS.n1315 DVSS.n758 4.06937
R9348 DVSS.n1321 DVSS.n758 4.06937
R9349 DVSS.n1321 DVSS.n627 4.06937
R9350 DVSS.n1337 DVSS.n627 4.06937
R9351 DVSS.n1337 DVSS.n628 4.06937
R9352 DVSS.n1333 DVSS.n628 4.06937
R9353 DVSS.n1333 DVSS.n1332 4.06937
R9354 DVSS.n1332 DVSS.n631 4.06937
R9355 DVSS.n662 DVSS.n631 4.06937
R9356 DVSS.n662 DVSS.n635 4.06937
R9357 DVSS.n753 DVSS.n635 4.06937
R9358 DVSS.n753 DVSS.n752 4.06937
R9359 DVSS.n752 DVSS.n638 4.06937
R9360 DVSS.n748 DVSS.n638 4.06937
R9361 DVSS.n748 DVSS.n747 4.06937
R9362 DVSS.n747 DVSS.n641 4.06937
R9363 DVSS.n743 DVSS.n641 4.06937
R9364 DVSS.n743 DVSS.n742 4.06937
R9365 DVSS.n742 DVSS.n644 4.06937
R9366 DVSS.n734 DVSS.n644 4.06937
R9367 DVSS.n734 DVSS.n733 4.06937
R9368 DVSS.n730 DVSS.n729 4.06937
R9369 DVSS.n729 DVSS.n650 4.06937
R9370 DVSS.n725 DVSS.n650 4.06937
R9371 DVSS.n725 DVSS.n724 4.06937
R9372 DVSS.n724 DVSS.n653 4.06937
R9373 DVSS.n720 DVSS.n653 4.06937
R9374 DVSS.n720 DVSS.n719 4.06937
R9375 DVSS.n719 DVSS.n656 4.06937
R9376 DVSS.n712 DVSS.n656 4.06937
R9377 DVSS.n712 DVSS.n711 4.06937
R9378 DVSS.n711 DVSS.n703 4.06937
R9379 DVSS.n703 DVSS.n541 4.06937
R9380 DVSS.n1657 DVSS.n541 4.06937
R9381 DVSS.n1657 DVSS.n539 4.06937
R9382 DVSS.n1666 DVSS.n539 4.06937
R9383 DVSS.n1666 DVSS.n536 4.06937
R9384 DVSS.n1672 DVSS.n536 4.06937
R9385 DVSS.n1672 DVSS.n535 4.06937
R9386 DVSS.n1677 DVSS.n535 4.06937
R9387 DVSS.n1677 DVSS.n531 4.06937
R9388 DVSS.n1684 DVSS.n531 4.06937
R9389 DVSS.n1684 DVSS.n530 4.06937
R9390 DVSS.n1694 DVSS.n530 4.06937
R9391 DVSS.n1694 DVSS.n527 4.06937
R9392 DVSS.n1700 DVSS.n527 4.06937
R9393 DVSS.n1705 DVSS.n526 4.06937
R9394 DVSS.n1705 DVSS.n522 4.06937
R9395 DVSS.n1712 DVSS.n522 4.06937
R9396 DVSS.n1712 DVSS.n521 4.06937
R9397 DVSS.n1717 DVSS.n521 4.06937
R9398 DVSS.n1717 DVSS.n513 4.06937
R9399 DVSS.n1739 DVSS.n513 4.06937
R9400 DVSS.n1739 DVSS.n1738 4.06937
R9401 DVSS.n1738 DVSS.n516 4.06937
R9402 DVSS.n1734 DVSS.n516 4.06937
R9403 DVSS.n1734 DVSS.n1733 4.06937
R9404 DVSS.n1733 DVSS.n509 4.06937
R9405 DVSS.n1750 DVSS.n509 4.06937
R9406 DVSS.n1750 DVSS.n505 4.06937
R9407 DVSS.n1757 DVSS.n505 4.06937
R9408 DVSS.n1757 DVSS.n504 4.06937
R9409 DVSS.n1762 DVSS.n504 4.06937
R9410 DVSS.n1762 DVSS.n500 4.06937
R9411 DVSS.n1768 DVSS.n500 4.06937
R9412 DVSS.n1768 DVSS.n499 4.06937
R9413 DVSS.n1773 DVSS.n499 4.06937
R9414 DVSS.n1773 DVSS.n495 4.06937
R9415 DVSS.n1781 DVSS.n495 4.06937
R9416 DVSS.n1788 DVSS.n1787 4.06937
R9417 DVSS.n1792 DVSS.n487 4.06937
R9418 DVSS.n1798 DVSS.n487 4.06937
R9419 DVSS.n1798 DVSS.n486 4.06937
R9420 DVSS.n1803 DVSS.n486 4.06937
R9421 DVSS.n1803 DVSS.n482 4.06937
R9422 DVSS.n1809 DVSS.n482 4.06937
R9423 DVSS.n1809 DVSS.n480 4.06937
R9424 DVSS.n1836 DVSS.n480 4.06937
R9425 DVSS.n1836 DVSS.n481 4.06937
R9426 DVSS.n1832 DVSS.n481 4.06937
R9427 DVSS.n1832 DVSS.n1831 4.06937
R9428 DVSS.n1831 DVSS.n1823 4.06937
R9429 DVSS.n1823 DVSS.n435 4.06937
R9430 DVSS.n1934 DVSS.n435 4.06937
R9431 DVSS.n1934 DVSS.n433 4.06937
R9432 DVSS.n1943 DVSS.n433 4.06937
R9433 DVSS.n1943 DVSS.n429 4.06937
R9434 DVSS.n1949 DVSS.n429 4.06937
R9435 DVSS.n1949 DVSS.n428 4.06937
R9436 DVSS.n1954 DVSS.n428 4.06937
R9437 DVSS.n1954 DVSS.n423 4.06937
R9438 DVSS.n1962 DVSS.n423 4.06937
R9439 DVSS.n1962 DVSS.n419 4.06937
R9440 DVSS.n1969 DVSS.n419 4.06937
R9441 DVSS.n1970 DVSS.n1969 4.06937
R9442 DVSS.n1974 DVSS.n415 4.06937
R9443 DVSS.n1980 DVSS.n415 4.06937
R9444 DVSS.n1980 DVSS.n414 4.06937
R9445 DVSS.n1985 DVSS.n414 4.06937
R9446 DVSS.n1985 DVSS.n410 4.06937
R9447 DVSS.n1991 DVSS.n410 4.06937
R9448 DVSS.n1991 DVSS.n408 4.06937
R9449 DVSS.n2018 DVSS.n408 4.06937
R9450 DVSS.n2018 DVSS.n409 4.06937
R9451 DVSS.n2014 DVSS.n409 4.06937
R9452 DVSS.n2014 DVSS.n2013 4.06937
R9453 DVSS.n2013 DVSS.n2005 4.06937
R9454 DVSS.n2005 DVSS.n363 4.06937
R9455 DVSS.n2116 DVSS.n363 4.06937
R9456 DVSS.n2116 DVSS.n361 4.06937
R9457 DVSS.n2125 DVSS.n361 4.06937
R9458 DVSS.n2125 DVSS.n357 4.06937
R9459 DVSS.n2131 DVSS.n357 4.06937
R9460 DVSS.n2131 DVSS.n356 4.06937
R9461 DVSS.n2136 DVSS.n356 4.06937
R9462 DVSS.n2136 DVSS.n351 4.06937
R9463 DVSS.n2144 DVSS.n351 4.06937
R9464 DVSS.n2144 DVSS.n347 4.06937
R9465 DVSS.n2151 DVSS.n347 4.06937
R9466 DVSS.n2152 DVSS.n2151 4.06937
R9467 DVSS.n2156 DVSS.n343 4.06937
R9468 DVSS.n2162 DVSS.n343 4.06937
R9469 DVSS.n2162 DVSS.n342 4.06937
R9470 DVSS.n2167 DVSS.n342 4.06937
R9471 DVSS.n2167 DVSS.n338 4.06937
R9472 DVSS.n2173 DVSS.n338 4.06937
R9473 DVSS.n2173 DVSS.n336 4.06937
R9474 DVSS.n2200 DVSS.n336 4.06937
R9475 DVSS.n2200 DVSS.n337 4.06937
R9476 DVSS.n2196 DVSS.n337 4.06937
R9477 DVSS.n2196 DVSS.n2195 4.06937
R9478 DVSS.n2195 DVSS.n2187 4.06937
R9479 DVSS.n2187 DVSS.n291 4.06937
R9480 DVSS.n2298 DVSS.n291 4.06937
R9481 DVSS.n2298 DVSS.n289 4.06937
R9482 DVSS.n2307 DVSS.n289 4.06937
R9483 DVSS.n2307 DVSS.n285 4.06937
R9484 DVSS.n2313 DVSS.n285 4.06937
R9485 DVSS.n2313 DVSS.n284 4.06937
R9486 DVSS.n2318 DVSS.n284 4.06937
R9487 DVSS.n2318 DVSS.n279 4.06937
R9488 DVSS.n2326 DVSS.n279 4.06937
R9489 DVSS.n2326 DVSS.n275 4.06937
R9490 DVSS.n2333 DVSS.n275 4.06937
R9491 DVSS.n2334 DVSS.n2333 4.06937
R9492 DVSS.n2338 DVSS.n271 4.06937
R9493 DVSS.n2344 DVSS.n271 4.06937
R9494 DVSS.n2344 DVSS.n270 4.06937
R9495 DVSS.n2349 DVSS.n270 4.06937
R9496 DVSS.n2349 DVSS.n266 4.06937
R9497 DVSS.n2355 DVSS.n266 4.06937
R9498 DVSS.n2355 DVSS.n135 4.06937
R9499 DVSS.n2371 DVSS.n135 4.06937
R9500 DVSS.n2371 DVSS.n136 4.06937
R9501 DVSS.n2367 DVSS.n136 4.06937
R9502 DVSS.n2367 DVSS.n2366 4.06937
R9503 DVSS.n2366 DVSS.n139 4.06937
R9504 DVSS.n170 DVSS.n139 4.06937
R9505 DVSS.n170 DVSS.n143 4.06937
R9506 DVSS.n261 DVSS.n143 4.06937
R9507 DVSS.n261 DVSS.n260 4.06937
R9508 DVSS.n260 DVSS.n146 4.06937
R9509 DVSS.n256 DVSS.n146 4.06937
R9510 DVSS.n256 DVSS.n255 4.06937
R9511 DVSS.n255 DVSS.n149 4.06937
R9512 DVSS.n251 DVSS.n149 4.06937
R9513 DVSS.n251 DVSS.n250 4.06937
R9514 DVSS.n250 DVSS.n152 4.06937
R9515 DVSS.n242 DVSS.n152 4.06937
R9516 DVSS.n242 DVSS.n241 4.06937
R9517 DVSS.n238 DVSS.n237 4.06937
R9518 DVSS.n237 DVSS.n158 4.06937
R9519 DVSS.n233 DVSS.n158 4.06937
R9520 DVSS.n233 DVSS.n232 4.06937
R9521 DVSS.n232 DVSS.n161 4.06937
R9522 DVSS.n228 DVSS.n161 4.06937
R9523 DVSS.n228 DVSS.n227 4.06937
R9524 DVSS.n227 DVSS.n164 4.06937
R9525 DVSS.n220 DVSS.n164 4.06937
R9526 DVSS.n220 DVSS.n219 4.06937
R9527 DVSS.n219 DVSS.n211 4.06937
R9528 DVSS.n211 DVSS.n49 4.06937
R9529 DVSS.n2650 DVSS.n49 4.06937
R9530 DVSS.n2650 DVSS.n47 4.06937
R9531 DVSS.n2659 DVSS.n47 4.06937
R9532 DVSS.n2659 DVSS.n44 4.06937
R9533 DVSS.n2665 DVSS.n44 4.06937
R9534 DVSS.n2665 DVSS.n43 4.06937
R9535 DVSS.n2670 DVSS.n43 4.06937
R9536 DVSS.n2670 DVSS.n39 4.06937
R9537 DVSS.n2677 DVSS.n39 4.06937
R9538 DVSS.n2677 DVSS.n38 4.06937
R9539 DVSS.n2687 DVSS.n38 4.06937
R9540 DVSS.n2687 DVSS.n35 4.06937
R9541 DVSS.n2693 DVSS.n35 4.06937
R9542 DVSS.n2698 DVSS.n34 4.06937
R9543 DVSS.n2698 DVSS.n30 4.06937
R9544 DVSS.n2705 DVSS.n30 4.06937
R9545 DVSS.n2705 DVSS.n29 4.06937
R9546 DVSS.n2710 DVSS.n29 4.06937
R9547 DVSS.n2710 DVSS.n21 4.06937
R9548 DVSS.n2732 DVSS.n21 4.06937
R9549 DVSS.n2732 DVSS.n2731 4.06937
R9550 DVSS.n2731 DVSS.n24 4.06937
R9551 DVSS.n2727 DVSS.n24 4.06937
R9552 DVSS.n2727 DVSS.n2726 4.06937
R9553 DVSS.n2726 DVSS.n17 4.06937
R9554 DVSS.n2743 DVSS.n17 4.06937
R9555 DVSS.n2743 DVSS.n13 4.06937
R9556 DVSS.n2750 DVSS.n13 4.06937
R9557 DVSS.n2750 DVSS.n11 4.06937
R9558 DVSS.n2781 DVSS.n11 4.06937
R9559 DVSS.n2781 DVSS.n12 4.06937
R9560 DVSS.n2777 DVSS.n12 4.06937
R9561 DVSS.n2777 DVSS.n2776 4.06937
R9562 DVSS.n2776 DVSS.n2755 4.06937
R9563 DVSS.n2772 DVSS.n2755 4.06937
R9564 DVSS.n2772 DVSS.n2771 4.06937
R9565 DVSS.n2771 DVSS.n2760 4.06937
R9566 DVSS.n2763 DVSS.n2760 4.06937
R9567 DVSS.n976 DVSS.n854 3.68864
R9568 DVSS.n1158 DVSS.n782 3.68864
R9569 DVSS.n1329 DVSS.n1326 3.68864
R9570 DVSS.n708 DVSS.n540 3.68864
R9571 DVSS.n1743 DVSS.n511 3.68864
R9572 DVSS.n1828 DVSS.n434 3.68864
R9573 DVSS.n2010 DVSS.n362 3.68864
R9574 DVSS.n2192 DVSS.n290 3.68864
R9575 DVSS.n2363 DVSS.n2360 3.68864
R9576 DVSS.n216 DVSS.n48 3.68864
R9577 DVSS.n2736 DVSS.n19 3.68864
R9578 DVSS.n1781 DVSS.n491 3.05216
R9579 DVSS.n1006 DVSS.n888 2.84494
R9580 DVSS.n1188 DVSS.n816 2.84494
R9581 DVSS.n1360 DVSS.n615 2.84494
R9582 DVSS.n1448 DVSS.n575 2.84494
R9583 DVSS.n1639 DVSS.n1638 2.84494
R9584 DVSS.n1858 DVSS.n468 2.84494
R9585 DVSS.n2040 DVSS.n396 2.84494
R9586 DVSS.n2222 DVSS.n324 2.84494
R9587 DVSS.n2394 DVSS.n123 2.84494
R9588 DVSS.n2482 DVSS.n83 2.84494
R9589 DVSS.n2632 DVSS.n2631 2.84494
R9590 DVSS.n888 DVSS 2.60791
R9591 DVSS.n816 DVSS 2.60791
R9592 DVSS.n615 DVSS 2.60791
R9593 DVSS.n575 DVSS 2.60791
R9594 DVSS.n1638 DVSS 2.60791
R9595 DVSS.n468 DVSS 2.60791
R9596 DVSS.n396 DVSS 2.60791
R9597 DVSS.n324 DVSS 2.60791
R9598 DVSS.n123 DVSS 2.60791
R9599 DVSS.n83 DVSS 2.60791
R9600 DVSS.n2631 DVSS 2.60791
R9601 DVSS.n934 DVSS.n913 2.38694
R9602 DVSS.n1057 DVSS.n868 2.38694
R9603 DVSS.n1239 DVSS.n796 2.38694
R9604 DVSS.n593 DVSS.n592 2.38694
R9605 DVSS.n1505 DVSS.n557 2.38694
R9606 DVSS.n1604 DVSS.n1603 2.38694
R9607 DVSS.n1909 DVSS.n448 2.38694
R9608 DVSS.n2091 DVSS.n376 2.38694
R9609 DVSS.n2273 DVSS.n304 2.38694
R9610 DVSS.n101 DVSS.n100 2.38694
R9611 DVSS.n2539 DVSS.n65 2.38694
R9612 DVSS.n1118 DVSS 2.03494
R9613 DVSS.n1122 DVSS 2.03494
R9614 DVSS.n1300 DVSS 2.03494
R9615 DVSS.n1304 DVSS 2.03494
R9616 DVSS.n733 DVSS 2.03494
R9617 DVSS.n730 DVSS 2.03494
R9618 DVSS.n1700 DVSS 2.03494
R9619 DVSS DVSS.n526 2.03494
R9620 DVSS.n1788 DVSS 2.03494
R9621 DVSS.n1792 DVSS 2.03494
R9622 DVSS.n1970 DVSS 2.03494
R9623 DVSS.n1974 DVSS 2.03494
R9624 DVSS.n2152 DVSS 2.03494
R9625 DVSS.n2156 DVSS 2.03494
R9626 DVSS.n2334 DVSS 2.03494
R9627 DVSS.n2338 DVSS 2.03494
R9628 DVSS.n241 DVSS 2.03494
R9629 DVSS.n238 DVSS 2.03494
R9630 DVSS.n2693 DVSS 2.03494
R9631 DVSS DVSS.n34 2.03494
R9632 DVSS.n2763 DVSS 2.03494
R9633 DVSS.n1039 DVSS 1.84457
R9634 DVSS DVSS.n1038 1.84457
R9635 DVSS.n1038 DVSS 1.84457
R9636 DVSS.n1221 DVSS 1.84457
R9637 DVSS DVSS.n1220 1.84457
R9638 DVSS.n1220 DVSS 1.84457
R9639 DVSS.n1396 DVSS 1.84457
R9640 DVSS DVSS.n1395 1.84457
R9641 DVSS.n1395 DVSS 1.84457
R9642 DVSS.n1483 DVSS 1.84457
R9643 DVSS DVSS.n1480 1.84457
R9644 DVSS.n1480 DVSS 1.84457
R9645 DVSS.n1616 DVSS 1.84457
R9646 DVSS DVSS.n1548 1.84457
R9647 DVSS.n1548 DVSS 1.84457
R9648 DVSS.n1891 DVSS 1.84457
R9649 DVSS DVSS.n1890 1.84457
R9650 DVSS.n1890 DVSS 1.84457
R9651 DVSS.n2073 DVSS 1.84457
R9652 DVSS DVSS.n2072 1.84457
R9653 DVSS.n2072 DVSS 1.84457
R9654 DVSS.n2255 DVSS 1.84457
R9655 DVSS DVSS.n2254 1.84457
R9656 DVSS.n2254 DVSS 1.84457
R9657 DVSS.n2430 DVSS 1.84457
R9658 DVSS DVSS.n2429 1.84457
R9659 DVSS.n2429 DVSS 1.84457
R9660 DVSS.n2517 DVSS 1.84457
R9661 DVSS DVSS.n2514 1.84457
R9662 DVSS.n2514 DVSS 1.84457
R9663 DVSS.n2609 DVSS 1.84457
R9664 DVSS DVSS.n2594 1.84457
R9665 DVSS.n2594 DVSS 1.84457
R9666 DVSS.n938 DVSS.n913 1.44683
R9667 DVSS.n1061 DVSS.n868 1.44683
R9668 DVSS.n1243 DVSS.n796 1.44683
R9669 DVSS.n592 DVSS.n591 1.44683
R9670 DVSS.n1509 DVSS.n557 1.44683
R9671 DVSS.n1603 DVSS.n1602 1.44683
R9672 DVSS.n1913 DVSS.n448 1.44683
R9673 DVSS.n2095 DVSS.n376 1.44683
R9674 DVSS.n2277 DVSS.n304 1.44683
R9675 DVSS.n100 DVSS.n99 1.44683
R9676 DVSS.n2543 DVSS.n65 1.44683
R9677 DVSS.n1025 DVSS.n877 1.34003
R9678 DVSS.n1037 DVSS.n877 1.34003
R9679 DVSS.n1023 DVSS.n883 1.34003
R9680 DVSS.n1207 DVSS.n805 1.34003
R9681 DVSS.n1219 DVSS.n805 1.34003
R9682 DVSS.n1205 DVSS.n811 1.34003
R9683 DVSS.n1379 DVSS.n605 1.34003
R9684 DVSS.n1394 DVSS.n605 1.34003
R9685 DVSS.n1377 DVSS.n610 1.34003
R9686 DVSS.n1465 DVSS.n566 1.34003
R9687 DVSS.n1479 DVSS.n566 1.34003
R9688 DVSS.n1463 DVSS.n570 1.34003
R9689 DVSS.n1624 DVSS.n1538 1.34003
R9690 DVSS.n1547 DVSS.n1538 1.34003
R9691 DVSS.n1626 DVSS.n1536 1.34003
R9692 DVSS.n1877 DVSS.n457 1.34003
R9693 DVSS.n1889 DVSS.n457 1.34003
R9694 DVSS.n1875 DVSS.n463 1.34003
R9695 DVSS.n2059 DVSS.n385 1.34003
R9696 DVSS.n2071 DVSS.n385 1.34003
R9697 DVSS.n2057 DVSS.n391 1.34003
R9698 DVSS.n2241 DVSS.n313 1.34003
R9699 DVSS.n2253 DVSS.n313 1.34003
R9700 DVSS.n2239 DVSS.n319 1.34003
R9701 DVSS.n2413 DVSS.n113 1.34003
R9702 DVSS.n2428 DVSS.n113 1.34003
R9703 DVSS.n2411 DVSS.n118 1.34003
R9704 DVSS.n2499 DVSS.n74 1.34003
R9705 DVSS.n2513 DVSS.n74 1.34003
R9706 DVSS.n2497 DVSS.n78 1.34003
R9707 DVSS.n2617 DVSS.n2580 1.34003
R9708 DVSS.n2593 DVSS.n2580 1.34003
R9709 DVSS.n2619 DVSS.n2578 1.34003
R9710 DVSS.n1778 DVSS.n491 1.3005
R9711 DVSS DVSS.n931 1.22087
R9712 DVSS.n1787 DVSS.n491 1.01772
R9713 DVSS.n933 DVSS 0.934277
R9714 DVSS.n1025 DVSS.n1024 0.856314
R9715 DVSS DVSS.n1037 0.856314
R9716 DVSS DVSS.n1023 0.856314
R9717 DVSS.n1207 DVSS.n1206 0.856314
R9718 DVSS DVSS.n1219 0.856314
R9719 DVSS DVSS.n1205 0.856314
R9720 DVSS.n1379 DVSS.n1378 0.856314
R9721 DVSS DVSS.n1394 0.856314
R9722 DVSS DVSS.n1377 0.856314
R9723 DVSS.n1465 DVSS.n1464 0.856314
R9724 DVSS DVSS.n1479 0.856314
R9725 DVSS DVSS.n1463 0.856314
R9726 DVSS.n1625 DVSS.n1624 0.856314
R9727 DVSS DVSS.n1547 0.856314
R9728 DVSS.n1626 DVSS 0.856314
R9729 DVSS.n1877 DVSS.n1876 0.856314
R9730 DVSS DVSS.n1889 0.856314
R9731 DVSS DVSS.n1875 0.856314
R9732 DVSS.n2059 DVSS.n2058 0.856314
R9733 DVSS DVSS.n2071 0.856314
R9734 DVSS DVSS.n2057 0.856314
R9735 DVSS.n2241 DVSS.n2240 0.856314
R9736 DVSS DVSS.n2253 0.856314
R9737 DVSS DVSS.n2239 0.856314
R9738 DVSS.n2413 DVSS.n2412 0.856314
R9739 DVSS DVSS.n2428 0.856314
R9740 DVSS DVSS.n2411 0.856314
R9741 DVSS.n2499 DVSS.n2498 0.856314
R9742 DVSS DVSS.n2513 0.856314
R9743 DVSS DVSS.n2497 0.856314
R9744 DVSS.n2618 DVSS.n2617 0.856314
R9745 DVSS DVSS.n2593 0.856314
R9746 DVSS.n2619 DVSS 0.856314
R9747 DVSS.n2762 DVSS 0.771333
R9748 DVSS.n2762 DVSS 0.479667
R9749 DVSS.n931 DVSS 0.110598
R9750 DVSS.n936 DVSS.n935 0.0714459
R9751 DVSS.n1059 DVSS.n1058 0.0714459
R9752 DVSS.n1241 DVSS.n1240 0.0714459
R9753 DVSS.n1414 DVSS.n594 0.0714459
R9754 DVSS.n1507 DVSS.n1506 0.0714459
R9755 DVSS.n1605 DVSS.n1557 0.0714459
R9756 DVSS.n1911 DVSS.n1910 0.0714459
R9757 DVSS.n2093 DVSS.n2092 0.0714459
R9758 DVSS.n2275 DVSS.n2274 0.0714459
R9759 DVSS.n2448 DVSS.n102 0.0714459
R9760 DVSS.n2541 DVSS.n2540 0.0714459
R9761 DVSS DVSS.n921 0.067223
R9762 DVSS.n958 DVSS 0.067223
R9763 DVSS.n959 DVSS 0.067223
R9764 DVSS DVSS.n982 0.067223
R9765 DVSS DVSS.n981 0.067223
R9766 DVSS DVSS.n972 0.067223
R9767 DVSS.n1090 DVSS 0.067223
R9768 DVSS DVSS.n1089 0.067223
R9769 DVSS.n1098 DVSS 0.067223
R9770 DVSS.n1099 DVSS 0.067223
R9771 DVSS.n1101 DVSS 0.067223
R9772 DVSS DVSS.n1100 0.067223
R9773 DVSS.n1111 DVSS 0.067223
R9774 DVSS.n1119 DVSS 0.067223
R9775 DVSS DVSS.n1131 0.067223
R9776 DVSS.n1140 DVSS 0.067223
R9777 DVSS.n1141 DVSS 0.067223
R9778 DVSS DVSS.n1164 0.067223
R9779 DVSS DVSS.n1163 0.067223
R9780 DVSS DVSS.n1154 0.067223
R9781 DVSS.n1272 DVSS 0.067223
R9782 DVSS DVSS.n1271 0.067223
R9783 DVSS.n1280 DVSS 0.067223
R9784 DVSS.n1281 DVSS 0.067223
R9785 DVSS.n1283 DVSS 0.067223
R9786 DVSS DVSS.n1282 0.067223
R9787 DVSS.n1293 DVSS 0.067223
R9788 DVSS.n1301 DVSS 0.067223
R9789 DVSS DVSS.n1313 0.067223
R9790 DVSS.n1322 DVSS 0.067223
R9791 DVSS.n1323 DVSS 0.067223
R9792 DVSS DVSS.n1335 0.067223
R9793 DVSS DVSS.n1334 0.067223
R9794 DVSS.n661 DVSS 0.067223
R9795 DVSS.n751 DVSS 0.067223
R9796 DVSS DVSS.n750 0.067223
R9797 DVSS DVSS.n749 0.067223
R9798 DVSS.n746 DVSS 0.067223
R9799 DVSS DVSS.n745 0.067223
R9800 DVSS DVSS.n744 0.067223
R9801 DVSS.n741 DVSS 0.067223
R9802 DVSS.n732 DVSS 0.067223
R9803 DVSS DVSS.n722 0.067223
R9804 DVSS DVSS.n721 0.067223
R9805 DVSS.n718 DVSS 0.067223
R9806 DVSS DVSS.n713 0.067223
R9807 DVSS.n710 DVSS 0.067223
R9808 DVSS.n1658 DVSS 0.067223
R9809 DVSS DVSS.n1664 0.067223
R9810 DVSS.n1673 DVSS 0.067223
R9811 DVSS.n1674 DVSS 0.067223
R9812 DVSS.n1676 DVSS 0.067223
R9813 DVSS DVSS.n1675 0.067223
R9814 DVSS.n1685 DVSS 0.067223
R9815 DVSS.n1686 DVSS 0.067223
R9816 DVSS.n1701 DVSS 0.067223
R9817 DVSS.n1716 DVSS 0.067223
R9818 DVSS DVSS.n1715 0.067223
R9819 DVSS.n1740 DVSS 0.067223
R9820 DVSS DVSS.n1736 0.067223
R9821 DVSS DVSS.n1735 0.067223
R9822 DVSS.n1749 DVSS 0.067223
R9823 DVSS.n1759 DVSS 0.067223
R9824 DVSS.n1761 DVSS 0.067223
R9825 DVSS DVSS.n1760 0.067223
R9826 DVSS.n1769 DVSS 0.067223
R9827 DVSS.n1770 DVSS 0.067223
R9828 DVSS.n1772 DVSS 0.067223
R9829 DVSS DVSS.n1771 0.067223
R9830 DVSS.n1789 DVSS 0.067223
R9831 DVSS DVSS.n1801 0.067223
R9832 DVSS.n1810 DVSS 0.067223
R9833 DVSS.n1811 DVSS 0.067223
R9834 DVSS DVSS.n1834 0.067223
R9835 DVSS DVSS.n1833 0.067223
R9836 DVSS DVSS.n1824 0.067223
R9837 DVSS.n1942 DVSS 0.067223
R9838 DVSS DVSS.n1941 0.067223
R9839 DVSS.n1950 DVSS 0.067223
R9840 DVSS.n1951 DVSS 0.067223
R9841 DVSS.n1953 DVSS 0.067223
R9842 DVSS DVSS.n1952 0.067223
R9843 DVSS.n1963 DVSS 0.067223
R9844 DVSS.n1971 DVSS 0.067223
R9845 DVSS DVSS.n1983 0.067223
R9846 DVSS.n1992 DVSS 0.067223
R9847 DVSS.n1993 DVSS 0.067223
R9848 DVSS DVSS.n2016 0.067223
R9849 DVSS DVSS.n2015 0.067223
R9850 DVSS DVSS.n2006 0.067223
R9851 DVSS.n2124 DVSS 0.067223
R9852 DVSS DVSS.n2123 0.067223
R9853 DVSS.n2132 DVSS 0.067223
R9854 DVSS.n2133 DVSS 0.067223
R9855 DVSS.n2135 DVSS 0.067223
R9856 DVSS DVSS.n2134 0.067223
R9857 DVSS.n2145 DVSS 0.067223
R9858 DVSS.n2153 DVSS 0.067223
R9859 DVSS DVSS.n2165 0.067223
R9860 DVSS.n2174 DVSS 0.067223
R9861 DVSS.n2175 DVSS 0.067223
R9862 DVSS DVSS.n2198 0.067223
R9863 DVSS DVSS.n2197 0.067223
R9864 DVSS DVSS.n2188 0.067223
R9865 DVSS.n2306 DVSS 0.067223
R9866 DVSS DVSS.n2305 0.067223
R9867 DVSS.n2314 DVSS 0.067223
R9868 DVSS.n2315 DVSS 0.067223
R9869 DVSS.n2317 DVSS 0.067223
R9870 DVSS DVSS.n2316 0.067223
R9871 DVSS.n2327 DVSS 0.067223
R9872 DVSS.n2335 DVSS 0.067223
R9873 DVSS DVSS.n2347 0.067223
R9874 DVSS.n2356 DVSS 0.067223
R9875 DVSS.n2357 DVSS 0.067223
R9876 DVSS DVSS.n2369 0.067223
R9877 DVSS DVSS.n2368 0.067223
R9878 DVSS.n169 DVSS 0.067223
R9879 DVSS.n259 DVSS 0.067223
R9880 DVSS DVSS.n258 0.067223
R9881 DVSS DVSS.n257 0.067223
R9882 DVSS.n254 DVSS 0.067223
R9883 DVSS DVSS.n253 0.067223
R9884 DVSS DVSS.n252 0.067223
R9885 DVSS.n249 DVSS 0.067223
R9886 DVSS.n240 DVSS 0.067223
R9887 DVSS DVSS.n230 0.067223
R9888 DVSS DVSS.n229 0.067223
R9889 DVSS.n226 DVSS 0.067223
R9890 DVSS DVSS.n221 0.067223
R9891 DVSS.n218 DVSS 0.067223
R9892 DVSS.n2651 DVSS 0.067223
R9893 DVSS DVSS.n2657 0.067223
R9894 DVSS.n2666 DVSS 0.067223
R9895 DVSS.n2667 DVSS 0.067223
R9896 DVSS.n2669 DVSS 0.067223
R9897 DVSS DVSS.n2668 0.067223
R9898 DVSS.n2678 DVSS 0.067223
R9899 DVSS.n2679 DVSS 0.067223
R9900 DVSS.n2694 DVSS 0.067223
R9901 DVSS.n2709 DVSS 0.067223
R9902 DVSS DVSS.n2708 0.067223
R9903 DVSS.n2733 DVSS 0.067223
R9904 DVSS DVSS.n2729 0.067223
R9905 DVSS DVSS.n2728 0.067223
R9906 DVSS.n2742 DVSS 0.067223
R9907 DVSS.n2752 DVSS 0.067223
R9908 DVSS.n2780 DVSS 0.067223
R9909 DVSS DVSS.n2779 0.067223
R9910 DVSS DVSS.n2778 0.067223
R9911 DVSS.n2775 DVSS 0.067223
R9912 DVSS DVSS.n2774 0.067223
R9913 DVSS DVSS.n2773 0.067223
R9914 DVSS DVSS.n2764 0.067223
R9915 DVSS.n942 DVSS.n909 0.067223
R9916 DVSS.n949 DVSS 0.067223
R9917 DVSS DVSS.n948 0.067223
R9918 DVSS.n992 DVSS 0.067223
R9919 DVSS.n993 DVSS 0.067223
R9920 DVSS.n995 DVSS 0.067223
R9921 DVSS DVSS.n994 0.067223
R9922 DVSS.n1012 DVSS 0.067223
R9923 DVSS DVSS.n1011 0.067223
R9924 DVSS.n1027 DVSS 0.067223
R9925 DVSS DVSS.n878 0.067223
R9926 DVSS.n1049 DVSS 0.067223
R9927 DVSS.n1050 DVSS 0.067223
R9928 DVSS.n1051 DVSS 0.067223
R9929 DVSS.n1065 DVSS.n864 0.067223
R9930 DVSS.n1072 DVSS 0.067223
R9931 DVSS DVSS.n1071 0.067223
R9932 DVSS.n1174 DVSS 0.067223
R9933 DVSS.n1175 DVSS 0.067223
R9934 DVSS.n1177 DVSS 0.067223
R9935 DVSS DVSS.n1176 0.067223
R9936 DVSS.n1194 DVSS 0.067223
R9937 DVSS DVSS.n1193 0.067223
R9938 DVSS.n1209 DVSS 0.067223
R9939 DVSS DVSS.n806 0.067223
R9940 DVSS.n1231 DVSS 0.067223
R9941 DVSS.n1232 DVSS 0.067223
R9942 DVSS.n1233 DVSS 0.067223
R9943 DVSS.n1247 DVSS.n792 0.067223
R9944 DVSS.n1254 DVSS 0.067223
R9945 DVSS DVSS.n1253 0.067223
R9946 DVSS.n1345 DVSS 0.067223
R9947 DVSS.n1346 DVSS 0.067223
R9948 DVSS.n1348 DVSS 0.067223
R9949 DVSS DVSS.n1347 0.067223
R9950 DVSS.n1366 DVSS 0.067223
R9951 DVSS DVSS.n1365 0.067223
R9952 DVSS.n1381 DVSS 0.067223
R9953 DVSS.n1389 DVSS 0.067223
R9954 DVSS DVSS.n1398 0.067223
R9955 DVSS.n1406 DVSS 0.067223
R9956 DVSS.n1407 DVSS 0.067223
R9957 DVSS.n1419 DVSS.n590 0.067223
R9958 DVSS DVSS.n1421 0.067223
R9959 DVSS.n1432 DVSS 0.067223
R9960 DVSS.n1433 DVSS 0.067223
R9961 DVSS.n1435 DVSS 0.067223
R9962 DVSS DVSS.n1434 0.067223
R9963 DVSS.n1444 DVSS 0.067223
R9964 DVSS DVSS.n1451 0.067223
R9965 DVSS.n1459 DVSS 0.067223
R9966 DVSS DVSS.n1467 0.067223
R9967 DVSS.n1485 DVSS 0.067223
R9968 DVSS.n1494 DVSS 0.067223
R9969 DVSS.n1496 DVSS 0.067223
R9970 DVSS DVSS.n1495 0.067223
R9971 DVSS.n1513 DVSS.n1512 0.067223
R9972 DVSS.n1522 DVSS 0.067223
R9973 DVSS.n1647 DVSS 0.067223
R9974 DVSS DVSS.n1646 0.067223
R9975 DVSS DVSS.n1645 0.067223
R9976 DVSS.n1642 DVSS 0.067223
R9977 DVSS DVSS.n1641 0.067223
R9978 DVSS DVSS.n1632 0.067223
R9979 DVSS DVSS.n1631 0.067223
R9980 DVSS.n1540 DVSS 0.067223
R9981 DVSS DVSS.n1618 0.067223
R9982 DVSS.n1611 DVSS 0.067223
R9983 DVSS DVSS.n1610 0.067223
R9984 DVSS DVSS.n1609 0.067223
R9985 DVSS.n1599 DVSS.n1560 0.067223
R9986 DVSS DVSS.n1594 0.067223
R9987 DVSS DVSS.n1564 0.067223
R9988 DVSS.n1844 DVSS 0.067223
R9989 DVSS.n1845 DVSS 0.067223
R9990 DVSS.n1847 DVSS 0.067223
R9991 DVSS DVSS.n1846 0.067223
R9992 DVSS.n1864 DVSS 0.067223
R9993 DVSS DVSS.n1863 0.067223
R9994 DVSS.n1879 DVSS 0.067223
R9995 DVSS DVSS.n458 0.067223
R9996 DVSS.n1901 DVSS 0.067223
R9997 DVSS.n1902 DVSS 0.067223
R9998 DVSS.n1903 DVSS 0.067223
R9999 DVSS.n1917 DVSS.n444 0.067223
R10000 DVSS.n1924 DVSS 0.067223
R10001 DVSS DVSS.n1923 0.067223
R10002 DVSS.n2026 DVSS 0.067223
R10003 DVSS.n2027 DVSS 0.067223
R10004 DVSS.n2029 DVSS 0.067223
R10005 DVSS DVSS.n2028 0.067223
R10006 DVSS.n2046 DVSS 0.067223
R10007 DVSS DVSS.n2045 0.067223
R10008 DVSS.n2061 DVSS 0.067223
R10009 DVSS DVSS.n386 0.067223
R10010 DVSS.n2083 DVSS 0.067223
R10011 DVSS.n2084 DVSS 0.067223
R10012 DVSS.n2085 DVSS 0.067223
R10013 DVSS.n2099 DVSS.n372 0.067223
R10014 DVSS.n2106 DVSS 0.067223
R10015 DVSS DVSS.n2105 0.067223
R10016 DVSS.n2208 DVSS 0.067223
R10017 DVSS.n2209 DVSS 0.067223
R10018 DVSS.n2211 DVSS 0.067223
R10019 DVSS DVSS.n2210 0.067223
R10020 DVSS.n2228 DVSS 0.067223
R10021 DVSS DVSS.n2227 0.067223
R10022 DVSS.n2243 DVSS 0.067223
R10023 DVSS DVSS.n314 0.067223
R10024 DVSS.n2265 DVSS 0.067223
R10025 DVSS.n2266 DVSS 0.067223
R10026 DVSS.n2267 DVSS 0.067223
R10027 DVSS.n2281 DVSS.n300 0.067223
R10028 DVSS.n2288 DVSS 0.067223
R10029 DVSS DVSS.n2287 0.067223
R10030 DVSS.n2379 DVSS 0.067223
R10031 DVSS.n2380 DVSS 0.067223
R10032 DVSS.n2382 DVSS 0.067223
R10033 DVSS DVSS.n2381 0.067223
R10034 DVSS.n2400 DVSS 0.067223
R10035 DVSS DVSS.n2399 0.067223
R10036 DVSS.n2415 DVSS 0.067223
R10037 DVSS.n2423 DVSS 0.067223
R10038 DVSS DVSS.n2432 0.067223
R10039 DVSS.n2440 DVSS 0.067223
R10040 DVSS.n2441 DVSS 0.067223
R10041 DVSS.n2453 DVSS.n98 0.067223
R10042 DVSS DVSS.n2455 0.067223
R10043 DVSS.n2466 DVSS 0.067223
R10044 DVSS.n2467 DVSS 0.067223
R10045 DVSS.n2469 DVSS 0.067223
R10046 DVSS DVSS.n2468 0.067223
R10047 DVSS.n2478 DVSS 0.067223
R10048 DVSS DVSS.n2485 0.067223
R10049 DVSS.n2493 DVSS 0.067223
R10050 DVSS DVSS.n2501 0.067223
R10051 DVSS.n2519 DVSS 0.067223
R10052 DVSS.n2528 DVSS 0.067223
R10053 DVSS.n2530 DVSS 0.067223
R10054 DVSS DVSS.n2529 0.067223
R10055 DVSS.n2547 DVSS.n2546 0.067223
R10056 DVSS.n2556 DVSS 0.067223
R10057 DVSS.n2640 DVSS 0.067223
R10058 DVSS DVSS.n2639 0.067223
R10059 DVSS DVSS.n2638 0.067223
R10060 DVSS.n2635 DVSS 0.067223
R10061 DVSS DVSS.n2634 0.067223
R10062 DVSS DVSS.n2625 0.067223
R10063 DVSS DVSS.n2624 0.067223
R10064 DVSS.n2582 DVSS 0.067223
R10065 DVSS DVSS.n2611 0.067223
R10066 DVSS.n2604 DVSS 0.067223
R10067 DVSS DVSS.n2603 0.067223
R10068 DVSS.n2787 DVSS 0.067223
R10069 DVSS DVSS.n1021 0.0663784
R10070 DVSS DVSS.n1203 0.0663784
R10071 DVSS DVSS.n1375 0.0663784
R10072 DVSS.n1468 DVSS 0.0663784
R10073 DVSS.n1539 DVSS 0.0663784
R10074 DVSS DVSS.n1873 0.0663784
R10075 DVSS DVSS.n2055 0.0663784
R10076 DVSS DVSS.n2237 0.0663784
R10077 DVSS DVSS.n2409 0.0663784
R10078 DVSS.n2502 DVSS 0.0663784
R10079 DVSS.n2581 DVSS 0.0663784
R10080 DVSS DVSS.n973 0.0638446
R10081 DVSS DVSS.n1155 0.0638446
R10082 DVSS.n660 DVSS 0.0638446
R10083 DVSS DVSS.n706 0.0638446
R10084 DVSS DVSS.n1730 0.0638446
R10085 DVSS DVSS.n1825 0.0638446
R10086 DVSS DVSS.n2007 0.0638446
R10087 DVSS DVSS.n2189 0.0638446
R10088 DVSS.n168 DVSS 0.0638446
R10089 DVSS DVSS.n214 0.0638446
R10090 DVSS DVSS.n2723 0.0638446
R10091 DVSS.n1113 DVSS 0.0613108
R10092 DVSS.n1295 DVSS 0.0613108
R10093 DVSS DVSS.n740 0.0613108
R10094 DVSS.n1687 DVSS 0.0613108
R10095 DVSS.n1783 DVSS 0.0613108
R10096 DVSS.n1965 DVSS 0.0613108
R10097 DVSS.n2147 DVSS 0.0613108
R10098 DVSS.n2329 DVSS 0.0613108
R10099 DVSS DVSS.n248 0.0613108
R10100 DVSS.n2680 DVSS 0.0613108
R10101 DVSS.n2761 DVSS 0.0613108
R10102 DVSS DVSS.n875 0.0477973
R10103 DVSS DVSS.n803 0.0477973
R10104 DVSS DVSS.n603 0.0477973
R10105 DVSS DVSS.n1484 0.0477973
R10106 DVSS DVSS.n1617 0.0477973
R10107 DVSS DVSS.n455 0.0477973
R10108 DVSS DVSS.n383 0.0477973
R10109 DVSS DVSS.n311 0.0477973
R10110 DVSS DVSS.n111 0.0477973
R10111 DVSS DVSS.n2518 0.0477973
R10112 DVSS DVSS.n2610 0.0477973
R10113 DVSS.n962 DVSS 0.0469527
R10114 DVSS.n1144 DVSS 0.0469527
R10115 DVSS DVSS.n757 0.0469527
R10116 DVSS.n715 DVSS 0.0469527
R10117 DVSS DVSS.n512 0.0469527
R10118 DVSS.n1814 DVSS 0.0469527
R10119 DVSS.n1996 DVSS 0.0469527
R10120 DVSS.n2178 DVSS 0.0469527
R10121 DVSS DVSS.n265 0.0469527
R10122 DVSS.n223 DVSS 0.0469527
R10123 DVSS DVSS.n20 0.0469527
R10124 DVSS DVSS.n1004 0.0469527
R10125 DVSS DVSS.n1186 0.0469527
R10126 DVSS DVSS.n1358 0.0469527
R10127 DVSS DVSS.n1446 0.0469527
R10128 DVSS.n1637 DVSS 0.0469527
R10129 DVSS DVSS.n1856 0.0469527
R10130 DVSS DVSS.n2038 0.0469527
R10131 DVSS DVSS.n2220 0.0469527
R10132 DVSS DVSS.n2392 0.0469527
R10133 DVSS DVSS.n2480 0.0469527
R10134 DVSS.n2630 DVSS 0.0469527
R10135 DVSS.n1020 DVSS 0.0461081
R10136 DVSS DVSS.n1035 0.0461081
R10137 DVSS.n1202 DVSS 0.0461081
R10138 DVSS DVSS.n1217 0.0461081
R10139 DVSS.n1374 DVSS 0.0461081
R10140 DVSS DVSS.n1392 0.0461081
R10141 DVSS.n1461 DVSS 0.0461081
R10142 DVSS DVSS.n1477 0.0461081
R10143 DVSS.n1628 DVSS 0.0461081
R10144 DVSS.n1619 DVSS 0.0461081
R10145 DVSS.n1872 DVSS 0.0461081
R10146 DVSS DVSS.n1887 0.0461081
R10147 DVSS.n2054 DVSS 0.0461081
R10148 DVSS DVSS.n2069 0.0461081
R10149 DVSS.n2236 DVSS 0.0461081
R10150 DVSS DVSS.n2251 0.0461081
R10151 DVSS.n2408 DVSS 0.0461081
R10152 DVSS DVSS.n2426 0.0461081
R10153 DVSS.n2495 DVSS 0.0461081
R10154 DVSS DVSS.n2511 0.0461081
R10155 DVSS.n2621 DVSS 0.0461081
R10156 DVSS.n2612 DVSS 0.0461081
R10157 DVSS.n978 DVSS 0.0435743
R10158 DVSS.n1088 DVSS 0.0435743
R10159 DVSS.n1160 DVSS 0.0435743
R10160 DVSS.n1270 DVSS 0.0435743
R10161 DVSS.n1331 DVSS 0.0435743
R10162 DVSS DVSS.n754 0.0435743
R10163 DVSS.n705 DVSS 0.0435743
R10164 DVSS.n1665 DVSS 0.0435743
R10165 DVSS.n1732 DVSS 0.0435743
R10166 DVSS.n1758 DVSS 0.0435743
R10167 DVSS.n1830 DVSS 0.0435743
R10168 DVSS.n1940 DVSS 0.0435743
R10169 DVSS.n2012 DVSS 0.0435743
R10170 DVSS.n2122 DVSS 0.0435743
R10171 DVSS.n2194 DVSS 0.0435743
R10172 DVSS.n2304 DVSS 0.0435743
R10173 DVSS.n2365 DVSS 0.0435743
R10174 DVSS DVSS.n262 0.0435743
R10175 DVSS.n213 DVSS 0.0435743
R10176 DVSS.n2658 DVSS 0.0435743
R10177 DVSS.n2725 DVSS 0.0435743
R10178 DVSS.n2751 DVSS 0.0435743
R10179 DVSS.n1008 DVSS 0.0418851
R10180 DVSS.n1190 DVSS 0.0418851
R10181 DVSS.n1362 DVSS 0.0418851
R10182 DVSS.n1450 DVSS 0.0418851
R10183 DVSS.n1531 DVSS 0.0418851
R10184 DVSS.n1860 DVSS 0.0418851
R10185 DVSS.n2042 DVSS 0.0418851
R10186 DVSS.n2224 DVSS 0.0418851
R10187 DVSS.n2396 DVSS 0.0418851
R10188 DVSS.n2484 DVSS 0.0418851
R10189 DVSS.n2571 DVSS 0.0418851
R10190 DVSS DVSS.n930 0.0410405
R10191 DVSS.n930 DVSS 0.0410405
R10192 DVSS.n919 DVSS 0.0410405
R10193 DVSS DVSS.n919 0.0410405
R10194 DVSS.n920 DVSS 0.0410405
R10195 DVSS DVSS.n920 0.0410405
R10196 DVSS.n922 DVSS 0.0410405
R10197 DVSS.n1115 DVSS 0.0410405
R10198 DVSS.n1121 DVSS 0.0410405
R10199 DVSS.n1121 DVSS 0.0410405
R10200 DVSS DVSS.n1120 0.0410405
R10201 DVSS.n1120 DVSS 0.0410405
R10202 DVSS.n1129 DVSS 0.0410405
R10203 DVSS DVSS.n1129 0.0410405
R10204 DVSS.n1130 DVSS 0.0410405
R10205 DVSS DVSS.n1130 0.0410405
R10206 DVSS.n1132 DVSS 0.0410405
R10207 DVSS.n1297 DVSS 0.0410405
R10208 DVSS.n1303 DVSS 0.0410405
R10209 DVSS.n1303 DVSS 0.0410405
R10210 DVSS DVSS.n1302 0.0410405
R10211 DVSS.n1302 DVSS 0.0410405
R10212 DVSS.n1311 DVSS 0.0410405
R10213 DVSS DVSS.n1311 0.0410405
R10214 DVSS.n1312 DVSS 0.0410405
R10215 DVSS DVSS.n1312 0.0410405
R10216 DVSS.n1314 DVSS 0.0410405
R10217 DVSS.n736 DVSS 0.0410405
R10218 DVSS DVSS.n731 0.0410405
R10219 DVSS.n731 DVSS 0.0410405
R10220 DVSS.n728 DVSS 0.0410405
R10221 DVSS.n728 DVSS 0.0410405
R10222 DVSS DVSS.n727 0.0410405
R10223 DVSS.n727 DVSS 0.0410405
R10224 DVSS DVSS.n726 0.0410405
R10225 DVSS.n726 DVSS 0.0410405
R10226 DVSS.n723 DVSS 0.0410405
R10227 DVSS DVSS.n1692 0.0410405
R10228 DVSS.n1702 DVSS 0.0410405
R10229 DVSS DVSS.n1702 0.0410405
R10230 DVSS.n1704 DVSS 0.0410405
R10231 DVSS.n1704 DVSS 0.0410405
R10232 DVSS DVSS.n1703 0.0410405
R10233 DVSS.n1703 DVSS 0.0410405
R10234 DVSS.n1713 DVSS 0.0410405
R10235 DVSS DVSS.n1713 0.0410405
R10236 DVSS.n1714 DVSS 0.0410405
R10237 DVSS.n1785 DVSS 0.0410405
R10238 DVSS.n1791 DVSS 0.0410405
R10239 DVSS.n1791 DVSS 0.0410405
R10240 DVSS DVSS.n1790 0.0410405
R10241 DVSS.n1790 DVSS 0.0410405
R10242 DVSS.n1799 DVSS 0.0410405
R10243 DVSS DVSS.n1799 0.0410405
R10244 DVSS.n1800 DVSS 0.0410405
R10245 DVSS DVSS.n1800 0.0410405
R10246 DVSS.n1802 DVSS 0.0410405
R10247 DVSS.n1967 DVSS 0.0410405
R10248 DVSS.n1973 DVSS 0.0410405
R10249 DVSS.n1973 DVSS 0.0410405
R10250 DVSS DVSS.n1972 0.0410405
R10251 DVSS.n1972 DVSS 0.0410405
R10252 DVSS.n1981 DVSS 0.0410405
R10253 DVSS DVSS.n1981 0.0410405
R10254 DVSS.n1982 DVSS 0.0410405
R10255 DVSS DVSS.n1982 0.0410405
R10256 DVSS.n1984 DVSS 0.0410405
R10257 DVSS.n2149 DVSS 0.0410405
R10258 DVSS.n2155 DVSS 0.0410405
R10259 DVSS.n2155 DVSS 0.0410405
R10260 DVSS DVSS.n2154 0.0410405
R10261 DVSS.n2154 DVSS 0.0410405
R10262 DVSS.n2163 DVSS 0.0410405
R10263 DVSS DVSS.n2163 0.0410405
R10264 DVSS.n2164 DVSS 0.0410405
R10265 DVSS DVSS.n2164 0.0410405
R10266 DVSS.n2166 DVSS 0.0410405
R10267 DVSS.n2331 DVSS 0.0410405
R10268 DVSS.n2337 DVSS 0.0410405
R10269 DVSS.n2337 DVSS 0.0410405
R10270 DVSS DVSS.n2336 0.0410405
R10271 DVSS.n2336 DVSS 0.0410405
R10272 DVSS.n2345 DVSS 0.0410405
R10273 DVSS DVSS.n2345 0.0410405
R10274 DVSS.n2346 DVSS 0.0410405
R10275 DVSS DVSS.n2346 0.0410405
R10276 DVSS.n2348 DVSS 0.0410405
R10277 DVSS.n244 DVSS 0.0410405
R10278 DVSS DVSS.n239 0.0410405
R10279 DVSS.n239 DVSS 0.0410405
R10280 DVSS.n236 DVSS 0.0410405
R10281 DVSS.n236 DVSS 0.0410405
R10282 DVSS DVSS.n235 0.0410405
R10283 DVSS.n235 DVSS 0.0410405
R10284 DVSS DVSS.n234 0.0410405
R10285 DVSS.n234 DVSS 0.0410405
R10286 DVSS.n231 DVSS 0.0410405
R10287 DVSS DVSS.n2685 0.0410405
R10288 DVSS.n2695 DVSS 0.0410405
R10289 DVSS DVSS.n2695 0.0410405
R10290 DVSS.n2697 DVSS 0.0410405
R10291 DVSS.n2697 DVSS 0.0410405
R10292 DVSS DVSS.n2696 0.0410405
R10293 DVSS.n2696 DVSS 0.0410405
R10294 DVSS.n2706 DVSS 0.0410405
R10295 DVSS DVSS.n2706 0.0410405
R10296 DVSS.n2707 DVSS 0.0410405
R10297 DVSS DVSS.n2769 0.0410405
R10298 DVSS DVSS.n946 0.0410405
R10299 DVSS.n947 DVSS 0.0410405
R10300 DVSS.n1056 DVSS 0.0410405
R10301 DVSS DVSS.n1069 0.0410405
R10302 DVSS.n1070 DVSS 0.0410405
R10303 DVSS.n1238 DVSS 0.0410405
R10304 DVSS DVSS.n1251 0.0410405
R10305 DVSS.n1252 DVSS 0.0410405
R10306 DVSS.n1408 DVSS 0.0410405
R10307 DVSS DVSS.n1420 0.0410405
R10308 DVSS.n1422 DVSS 0.0410405
R10309 DVSS.n1504 DVSS 0.0410405
R10310 DVSS.n556 DVSS 0.0410405
R10311 DVSS.n1521 DVSS 0.0410405
R10312 DVSS.n1606 DVSS 0.0410405
R10313 DVSS.n1596 DVSS 0.0410405
R10314 DVSS DVSS.n1595 0.0410405
R10315 DVSS.n1908 DVSS 0.0410405
R10316 DVSS DVSS.n1921 0.0410405
R10317 DVSS.n1922 DVSS 0.0410405
R10318 DVSS.n2090 DVSS 0.0410405
R10319 DVSS DVSS.n2103 0.0410405
R10320 DVSS.n2104 DVSS 0.0410405
R10321 DVSS.n2272 DVSS 0.0410405
R10322 DVSS DVSS.n2285 0.0410405
R10323 DVSS.n2286 DVSS 0.0410405
R10324 DVSS.n2442 DVSS 0.0410405
R10325 DVSS DVSS.n2454 0.0410405
R10326 DVSS.n2456 DVSS 0.0410405
R10327 DVSS.n2538 DVSS 0.0410405
R10328 DVSS.n64 DVSS 0.0410405
R10329 DVSS.n2555 DVSS 0.0410405
R10330 DVSS.n937 DVSS 0.0376622
R10331 DVSS.n941 DVSS 0.0376622
R10332 DVSS.n1060 DVSS 0.0376622
R10333 DVSS.n1064 DVSS 0.0376622
R10334 DVSS.n1242 DVSS 0.0376622
R10335 DVSS.n1246 DVSS 0.0376622
R10336 DVSS DVSS.n1415 0.0376622
R10337 DVSS.n1416 DVSS 0.0376622
R10338 DVSS.n1508 DVSS 0.0376622
R10339 DVSS DVSS.n555 0.0376622
R10340 DVSS.n1601 DVSS 0.0376622
R10341 DVSS DVSS.n1600 0.0376622
R10342 DVSS.n1912 DVSS 0.0376622
R10343 DVSS.n1916 DVSS 0.0376622
R10344 DVSS.n2094 DVSS 0.0376622
R10345 DVSS.n2098 DVSS 0.0376622
R10346 DVSS.n2276 DVSS 0.0376622
R10347 DVSS.n2280 DVSS 0.0376622
R10348 DVSS DVSS.n2449 0.0376622
R10349 DVSS.n2450 DVSS 0.0376622
R10350 DVSS.n2542 DVSS 0.0376622
R10351 DVSS DVSS.n63 0.0376622
R10352 DVSS.n1084 DVSS 0.0300608
R10353 DVSS.n1266 DVSS 0.0300608
R10354 DVSS DVSS.n632 0.0300608
R10355 DVSS.n1660 DVSS 0.0300608
R10356 DVSS DVSS.n1748 0.0300608
R10357 DVSS.n1936 DVSS 0.0300608
R10358 DVSS.n2118 DVSS 0.0300608
R10359 DVSS.n2300 DVSS 0.0300608
R10360 DVSS DVSS.n140 0.0300608
R10361 DVSS.n2653 DVSS 0.0300608
R10362 DVSS DVSS.n2741 0.0300608
R10363 DVSS DVSS.n1026 0.027527
R10364 DVSS DVSS.n1040 0.027527
R10365 DVSS DVSS.n1208 0.027527
R10366 DVSS DVSS.n1222 0.027527
R10367 DVSS DVSS.n1380 0.027527
R10368 DVSS.n1397 DVSS 0.027527
R10369 DVSS DVSS.n1466 0.027527
R10370 DVSS.n1482 DVSS 0.027527
R10371 DVSS.n1623 DVSS 0.027527
R10372 DVSS.n1615 DVSS 0.027527
R10373 DVSS DVSS.n1878 0.027527
R10374 DVSS DVSS.n1892 0.027527
R10375 DVSS DVSS.n2060 0.027527
R10376 DVSS DVSS.n2074 0.027527
R10377 DVSS DVSS.n2242 0.027527
R10378 DVSS DVSS.n2256 0.027527
R10379 DVSS DVSS.n2414 0.027527
R10380 DVSS.n2431 DVSS 0.027527
R10381 DVSS DVSS.n2500 0.027527
R10382 DVSS.n2516 DVSS 0.027527
R10383 DVSS.n2616 DVSS 0.027527
R10384 DVSS.n2608 DVSS 0.027527
R10385 DVSS DVSS.n882 0.0258378
R10386 DVSS DVSS.n873 0.0258378
R10387 DVSS DVSS.n810 0.0258378
R10388 DVSS DVSS.n801 0.0258378
R10389 DVSS DVSS.n609 0.0258378
R10390 DVSS.n1399 DVSS 0.0258378
R10391 DVSS.n1476 DVSS 0.0258378
R10392 DVSS.n1493 DVSS 0.0258378
R10393 DVSS DVSS.n1622 0.0258378
R10394 DVSS DVSS.n1614 0.0258378
R10395 DVSS DVSS.n462 0.0258378
R10396 DVSS DVSS.n453 0.0258378
R10397 DVSS DVSS.n390 0.0258378
R10398 DVSS DVSS.n381 0.0258378
R10399 DVSS DVSS.n318 0.0258378
R10400 DVSS DVSS.n309 0.0258378
R10401 DVSS DVSS.n117 0.0258378
R10402 DVSS.n2433 DVSS 0.0258378
R10403 DVSS.n2510 DVSS 0.0258378
R10404 DVSS.n2527 DVSS 0.0258378
R10405 DVSS DVSS.n2615 0.0258378
R10406 DVSS DVSS.n2607 0.0258378
R10407 DVSS DVSS.n1083 0.0233041
R10408 DVSS DVSS.n1265 0.0233041
R10409 DVSS.n634 DVSS 0.0233041
R10410 DVSS DVSS.n1659 0.0233041
R10411 DVSS.n1745 DVSS 0.0233041
R10412 DVSS DVSS.n1935 0.0233041
R10413 DVSS DVSS.n2117 0.0233041
R10414 DVSS DVSS.n2299 0.0233041
R10415 DVSS.n142 DVSS 0.0233041
R10416 DVSS DVSS.n2652 0.0233041
R10417 DVSS.n2738 DVSS 0.0233041
R10418 DVSS DVSS.n2762 0.0216149
R10419 DVSS.n922 DVSS 0.0148581
R10420 DVSS.n921 DVSS 0.0148581
R10421 DVSS DVSS.n958 0.0148581
R10422 DVSS DVSS.n962 0.0148581
R10423 DVSS.n983 DVSS 0.0148581
R10424 DVSS.n982 DVSS 0.0148581
R10425 DVSS.n981 DVSS 0.0148581
R10426 DVSS.n974 DVSS 0.0148581
R10427 DVSS.n973 DVSS 0.0148581
R10428 DVSS.n972 DVSS 0.0148581
R10429 DVSS.n1084 DVSS 0.0148581
R10430 DVSS.n1083 DVSS 0.0148581
R10431 DVSS DVSS.n1087 0.0148581
R10432 DVSS DVSS.n1088 0.0148581
R10433 DVSS.n1090 DVSS 0.0148581
R10434 DVSS.n1089 DVSS 0.0148581
R10435 DVSS DVSS.n1098 0.0148581
R10436 DVSS DVSS.n1099 0.0148581
R10437 DVSS.n1101 DVSS 0.0148581
R10438 DVSS.n1100 DVSS 0.0148581
R10439 DVSS DVSS.n1111 0.0148581
R10440 DVSS DVSS.n1115 0.0148581
R10441 DVSS.n1116 DVSS 0.0148581
R10442 DVSS DVSS.n1119 0.0148581
R10443 DVSS.n1132 DVSS 0.0148581
R10444 DVSS.n1131 DVSS 0.0148581
R10445 DVSS DVSS.n1140 0.0148581
R10446 DVSS DVSS.n1144 0.0148581
R10447 DVSS.n1165 DVSS 0.0148581
R10448 DVSS.n1164 DVSS 0.0148581
R10449 DVSS.n1163 DVSS 0.0148581
R10450 DVSS.n1156 DVSS 0.0148581
R10451 DVSS.n1155 DVSS 0.0148581
R10452 DVSS.n1154 DVSS 0.0148581
R10453 DVSS.n1266 DVSS 0.0148581
R10454 DVSS.n1265 DVSS 0.0148581
R10455 DVSS DVSS.n1269 0.0148581
R10456 DVSS DVSS.n1270 0.0148581
R10457 DVSS.n1272 DVSS 0.0148581
R10458 DVSS.n1271 DVSS 0.0148581
R10459 DVSS DVSS.n1280 0.0148581
R10460 DVSS DVSS.n1281 0.0148581
R10461 DVSS.n1283 DVSS 0.0148581
R10462 DVSS.n1282 DVSS 0.0148581
R10463 DVSS DVSS.n1293 0.0148581
R10464 DVSS DVSS.n1297 0.0148581
R10465 DVSS.n1298 DVSS 0.0148581
R10466 DVSS DVSS.n1301 0.0148581
R10467 DVSS.n1314 DVSS 0.0148581
R10468 DVSS.n1313 DVSS 0.0148581
R10469 DVSS DVSS.n1322 0.0148581
R10470 DVSS.n757 DVSS 0.0148581
R10471 DVSS.n1336 DVSS 0.0148581
R10472 DVSS.n1335 DVSS 0.0148581
R10473 DVSS.n1334 DVSS 0.0148581
R10474 DVSS.n1327 DVSS 0.0148581
R10475 DVSS DVSS.n660 0.0148581
R10476 DVSS.n661 DVSS 0.0148581
R10477 DVSS DVSS.n632 0.0148581
R10478 DVSS.n634 DVSS 0.0148581
R10479 DVSS.n755 DVSS 0.0148581
R10480 DVSS.n754 DVSS 0.0148581
R10481 DVSS.n751 DVSS 0.0148581
R10482 DVSS.n750 DVSS 0.0148581
R10483 DVSS.n749 DVSS 0.0148581
R10484 DVSS.n746 DVSS 0.0148581
R10485 DVSS.n745 DVSS 0.0148581
R10486 DVSS.n744 DVSS 0.0148581
R10487 DVSS.n741 DVSS 0.0148581
R10488 DVSS.n736 DVSS 0.0148581
R10489 DVSS.n735 DVSS 0.0148581
R10490 DVSS.n732 DVSS 0.0148581
R10491 DVSS.n723 DVSS 0.0148581
R10492 DVSS.n722 DVSS 0.0148581
R10493 DVSS.n721 DVSS 0.0148581
R10494 DVSS.n715 DVSS 0.0148581
R10495 DVSS.n714 DVSS 0.0148581
R10496 DVSS.n713 DVSS 0.0148581
R10497 DVSS.n710 DVSS 0.0148581
R10498 DVSS.n709 DVSS 0.0148581
R10499 DVSS.n706 DVSS 0.0148581
R10500 DVSS DVSS.n1658 0.0148581
R10501 DVSS.n1660 DVSS 0.0148581
R10502 DVSS.n1659 DVSS 0.0148581
R10503 DVSS DVSS.n1663 0.0148581
R10504 DVSS.n1665 DVSS 0.0148581
R10505 DVSS.n1664 DVSS 0.0148581
R10506 DVSS DVSS.n1673 0.0148581
R10507 DVSS DVSS.n1674 0.0148581
R10508 DVSS.n1676 DVSS 0.0148581
R10509 DVSS.n1675 DVSS 0.0148581
R10510 DVSS DVSS.n1685 0.0148581
R10511 DVSS DVSS.n1686 0.0148581
R10512 DVSS.n1692 DVSS 0.0148581
R10513 DVSS.n1688 DVSS 0.0148581
R10514 DVSS DVSS.n1701 0.0148581
R10515 DVSS DVSS.n1714 0.0148581
R10516 DVSS.n1716 DVSS 0.0148581
R10517 DVSS.n1715 DVSS 0.0148581
R10518 DVSS DVSS.n512 0.0148581
R10519 DVSS.n1737 DVSS 0.0148581
R10520 DVSS.n1736 DVSS 0.0148581
R10521 DVSS.n1735 DVSS 0.0148581
R10522 DVSS DVSS.n1729 0.0148581
R10523 DVSS.n1730 DVSS 0.0148581
R10524 DVSS.n1749 DVSS 0.0148581
R10525 DVSS.n1748 DVSS 0.0148581
R10526 DVSS DVSS.n1745 0.0148581
R10527 DVSS.n1746 DVSS 0.0148581
R10528 DVSS DVSS.n1758 0.0148581
R10529 DVSS DVSS.n1759 0.0148581
R10530 DVSS.n1761 DVSS 0.0148581
R10531 DVSS.n1760 DVSS 0.0148581
R10532 DVSS DVSS.n1769 0.0148581
R10533 DVSS DVSS.n1770 0.0148581
R10534 DVSS.n1772 DVSS 0.0148581
R10535 DVSS.n1771 DVSS 0.0148581
R10536 DVSS DVSS.n1785 0.0148581
R10537 DVSS.n1786 DVSS 0.0148581
R10538 DVSS DVSS.n1789 0.0148581
R10539 DVSS.n1802 DVSS 0.0148581
R10540 DVSS.n1801 DVSS 0.0148581
R10541 DVSS DVSS.n1810 0.0148581
R10542 DVSS DVSS.n1814 0.0148581
R10543 DVSS.n1835 DVSS 0.0148581
R10544 DVSS.n1834 DVSS 0.0148581
R10545 DVSS.n1833 DVSS 0.0148581
R10546 DVSS.n1826 DVSS 0.0148581
R10547 DVSS.n1825 DVSS 0.0148581
R10548 DVSS.n1824 DVSS 0.0148581
R10549 DVSS.n1936 DVSS 0.0148581
R10550 DVSS.n1935 DVSS 0.0148581
R10551 DVSS DVSS.n1939 0.0148581
R10552 DVSS DVSS.n1940 0.0148581
R10553 DVSS.n1942 DVSS 0.0148581
R10554 DVSS.n1941 DVSS 0.0148581
R10555 DVSS DVSS.n1950 0.0148581
R10556 DVSS DVSS.n1951 0.0148581
R10557 DVSS.n1953 DVSS 0.0148581
R10558 DVSS.n1952 DVSS 0.0148581
R10559 DVSS DVSS.n1963 0.0148581
R10560 DVSS DVSS.n1967 0.0148581
R10561 DVSS.n1968 DVSS 0.0148581
R10562 DVSS DVSS.n1971 0.0148581
R10563 DVSS.n1984 DVSS 0.0148581
R10564 DVSS.n1983 DVSS 0.0148581
R10565 DVSS DVSS.n1992 0.0148581
R10566 DVSS DVSS.n1996 0.0148581
R10567 DVSS.n2017 DVSS 0.0148581
R10568 DVSS.n2016 DVSS 0.0148581
R10569 DVSS.n2015 DVSS 0.0148581
R10570 DVSS.n2008 DVSS 0.0148581
R10571 DVSS.n2007 DVSS 0.0148581
R10572 DVSS.n2006 DVSS 0.0148581
R10573 DVSS.n2118 DVSS 0.0148581
R10574 DVSS.n2117 DVSS 0.0148581
R10575 DVSS DVSS.n2121 0.0148581
R10576 DVSS DVSS.n2122 0.0148581
R10577 DVSS.n2124 DVSS 0.0148581
R10578 DVSS.n2123 DVSS 0.0148581
R10579 DVSS DVSS.n2132 0.0148581
R10580 DVSS DVSS.n2133 0.0148581
R10581 DVSS.n2135 DVSS 0.0148581
R10582 DVSS.n2134 DVSS 0.0148581
R10583 DVSS DVSS.n2145 0.0148581
R10584 DVSS DVSS.n2149 0.0148581
R10585 DVSS.n2150 DVSS 0.0148581
R10586 DVSS DVSS.n2153 0.0148581
R10587 DVSS.n2166 DVSS 0.0148581
R10588 DVSS.n2165 DVSS 0.0148581
R10589 DVSS DVSS.n2174 0.0148581
R10590 DVSS DVSS.n2178 0.0148581
R10591 DVSS.n2199 DVSS 0.0148581
R10592 DVSS.n2198 DVSS 0.0148581
R10593 DVSS.n2197 DVSS 0.0148581
R10594 DVSS.n2190 DVSS 0.0148581
R10595 DVSS.n2189 DVSS 0.0148581
R10596 DVSS.n2188 DVSS 0.0148581
R10597 DVSS.n2300 DVSS 0.0148581
R10598 DVSS.n2299 DVSS 0.0148581
R10599 DVSS DVSS.n2303 0.0148581
R10600 DVSS DVSS.n2304 0.0148581
R10601 DVSS.n2306 DVSS 0.0148581
R10602 DVSS.n2305 DVSS 0.0148581
R10603 DVSS DVSS.n2314 0.0148581
R10604 DVSS DVSS.n2315 0.0148581
R10605 DVSS.n2317 DVSS 0.0148581
R10606 DVSS.n2316 DVSS 0.0148581
R10607 DVSS DVSS.n2327 0.0148581
R10608 DVSS DVSS.n2331 0.0148581
R10609 DVSS.n2332 DVSS 0.0148581
R10610 DVSS DVSS.n2335 0.0148581
R10611 DVSS.n2348 DVSS 0.0148581
R10612 DVSS.n2347 DVSS 0.0148581
R10613 DVSS DVSS.n2356 0.0148581
R10614 DVSS.n265 DVSS 0.0148581
R10615 DVSS.n2370 DVSS 0.0148581
R10616 DVSS.n2369 DVSS 0.0148581
R10617 DVSS.n2368 DVSS 0.0148581
R10618 DVSS.n2361 DVSS 0.0148581
R10619 DVSS DVSS.n168 0.0148581
R10620 DVSS.n169 DVSS 0.0148581
R10621 DVSS DVSS.n140 0.0148581
R10622 DVSS.n142 DVSS 0.0148581
R10623 DVSS.n263 DVSS 0.0148581
R10624 DVSS.n262 DVSS 0.0148581
R10625 DVSS.n259 DVSS 0.0148581
R10626 DVSS.n258 DVSS 0.0148581
R10627 DVSS.n257 DVSS 0.0148581
R10628 DVSS.n254 DVSS 0.0148581
R10629 DVSS.n253 DVSS 0.0148581
R10630 DVSS.n252 DVSS 0.0148581
R10631 DVSS.n249 DVSS 0.0148581
R10632 DVSS.n244 DVSS 0.0148581
R10633 DVSS.n243 DVSS 0.0148581
R10634 DVSS.n240 DVSS 0.0148581
R10635 DVSS.n231 DVSS 0.0148581
R10636 DVSS.n230 DVSS 0.0148581
R10637 DVSS.n229 DVSS 0.0148581
R10638 DVSS.n223 DVSS 0.0148581
R10639 DVSS.n222 DVSS 0.0148581
R10640 DVSS.n221 DVSS 0.0148581
R10641 DVSS.n218 DVSS 0.0148581
R10642 DVSS.n217 DVSS 0.0148581
R10643 DVSS.n214 DVSS 0.0148581
R10644 DVSS DVSS.n2651 0.0148581
R10645 DVSS.n2653 DVSS 0.0148581
R10646 DVSS.n2652 DVSS 0.0148581
R10647 DVSS DVSS.n2656 0.0148581
R10648 DVSS.n2658 DVSS 0.0148581
R10649 DVSS.n2657 DVSS 0.0148581
R10650 DVSS DVSS.n2666 0.0148581
R10651 DVSS DVSS.n2667 0.0148581
R10652 DVSS.n2669 DVSS 0.0148581
R10653 DVSS.n2668 DVSS 0.0148581
R10654 DVSS DVSS.n2678 0.0148581
R10655 DVSS DVSS.n2679 0.0148581
R10656 DVSS.n2685 DVSS 0.0148581
R10657 DVSS.n2681 DVSS 0.0148581
R10658 DVSS DVSS.n2694 0.0148581
R10659 DVSS DVSS.n2707 0.0148581
R10660 DVSS.n2709 DVSS 0.0148581
R10661 DVSS.n2708 DVSS 0.0148581
R10662 DVSS DVSS.n20 0.0148581
R10663 DVSS.n2730 DVSS 0.0148581
R10664 DVSS.n2729 DVSS 0.0148581
R10665 DVSS.n2728 DVSS 0.0148581
R10666 DVSS DVSS.n2722 0.0148581
R10667 DVSS.n2723 DVSS 0.0148581
R10668 DVSS.n2742 DVSS 0.0148581
R10669 DVSS.n2741 DVSS 0.0148581
R10670 DVSS DVSS.n2738 0.0148581
R10671 DVSS.n2739 DVSS 0.0148581
R10672 DVSS DVSS.n2751 0.0148581
R10673 DVSS DVSS.n2752 0.0148581
R10674 DVSS.n2780 DVSS 0.0148581
R10675 DVSS.n2779 DVSS 0.0148581
R10676 DVSS.n2778 DVSS 0.0148581
R10677 DVSS.n2775 DVSS 0.0148581
R10678 DVSS.n2774 DVSS 0.0148581
R10679 DVSS.n2773 DVSS 0.0148581
R10680 DVSS.n2769 DVSS 0.0148581
R10681 DVSS.n2765 DVSS 0.0148581
R10682 DVSS.n2764 DVSS 0.0148581
R10683 DVSS.n946 DVSS.n909 0.0148581
R10684 DVSS DVSS.n947 0.0148581
R10685 DVSS.n949 DVSS 0.0148581
R10686 DVSS.n948 DVSS 0.0148581
R10687 DVSS DVSS.n992 0.0148581
R10688 DVSS DVSS.n993 0.0148581
R10689 DVSS.n995 DVSS 0.0148581
R10690 DVSS.n994 DVSS 0.0148581
R10691 DVSS.n1005 DVSS 0.0148581
R10692 DVSS DVSS.n1008 0.0148581
R10693 DVSS DVSS.n1009 0.0148581
R10694 DVSS.n1012 DVSS 0.0148581
R10695 DVSS.n1011 DVSS 0.0148581
R10696 DVSS.n1010 DVSS 0.0148581
R10697 DVSS.n1021 DVSS 0.0148581
R10698 DVSS.n1027 DVSS 0.0148581
R10699 DVSS.n1026 DVSS 0.0148581
R10700 DVSS.n882 DVSS 0.0148581
R10701 DVSS.n1036 DVSS 0.0148581
R10702 DVSS.n1035 DVSS 0.0148581
R10703 DVSS.n878 DVSS 0.0148581
R10704 DVSS.n875 DVSS 0.0148581
R10705 DVSS.n1041 DVSS 0.0148581
R10706 DVSS.n1040 DVSS 0.0148581
R10707 DVSS.n873 DVSS 0.0148581
R10708 DVSS DVSS.n1049 0.0148581
R10709 DVSS DVSS.n1050 0.0148581
R10710 DVSS.n1051 DVSS 0.0148581
R10711 DVSS.n1069 DVSS.n864 0.0148581
R10712 DVSS DVSS.n1070 0.0148581
R10713 DVSS.n1072 DVSS 0.0148581
R10714 DVSS.n1071 DVSS 0.0148581
R10715 DVSS DVSS.n1174 0.0148581
R10716 DVSS DVSS.n1175 0.0148581
R10717 DVSS.n1177 DVSS 0.0148581
R10718 DVSS.n1176 DVSS 0.0148581
R10719 DVSS.n1187 DVSS 0.0148581
R10720 DVSS DVSS.n1190 0.0148581
R10721 DVSS DVSS.n1191 0.0148581
R10722 DVSS.n1194 DVSS 0.0148581
R10723 DVSS.n1193 DVSS 0.0148581
R10724 DVSS.n1192 DVSS 0.0148581
R10725 DVSS.n1203 DVSS 0.0148581
R10726 DVSS.n1209 DVSS 0.0148581
R10727 DVSS.n1208 DVSS 0.0148581
R10728 DVSS.n810 DVSS 0.0148581
R10729 DVSS.n1218 DVSS 0.0148581
R10730 DVSS.n1217 DVSS 0.0148581
R10731 DVSS.n806 DVSS 0.0148581
R10732 DVSS.n803 DVSS 0.0148581
R10733 DVSS.n1223 DVSS 0.0148581
R10734 DVSS.n1222 DVSS 0.0148581
R10735 DVSS.n801 DVSS 0.0148581
R10736 DVSS DVSS.n1231 0.0148581
R10737 DVSS DVSS.n1232 0.0148581
R10738 DVSS.n1233 DVSS 0.0148581
R10739 DVSS.n1251 DVSS.n792 0.0148581
R10740 DVSS DVSS.n1252 0.0148581
R10741 DVSS.n1254 DVSS 0.0148581
R10742 DVSS.n1253 DVSS 0.0148581
R10743 DVSS DVSS.n1345 0.0148581
R10744 DVSS DVSS.n1346 0.0148581
R10745 DVSS.n1348 DVSS 0.0148581
R10746 DVSS.n1347 DVSS 0.0148581
R10747 DVSS.n1359 DVSS 0.0148581
R10748 DVSS DVSS.n1362 0.0148581
R10749 DVSS DVSS.n1363 0.0148581
R10750 DVSS.n1366 DVSS 0.0148581
R10751 DVSS.n1365 DVSS 0.0148581
R10752 DVSS.n1364 DVSS 0.0148581
R10753 DVSS.n1375 DVSS 0.0148581
R10754 DVSS.n1381 DVSS 0.0148581
R10755 DVSS.n1380 DVSS 0.0148581
R10756 DVSS.n609 DVSS 0.0148581
R10757 DVSS.n1393 DVSS 0.0148581
R10758 DVSS.n1392 DVSS 0.0148581
R10759 DVSS.n1389 DVSS 0.0148581
R10760 DVSS.n603 DVSS 0.0148581
R10761 DVSS.n602 DVSS 0.0148581
R10762 DVSS DVSS.n1397 0.0148581
R10763 DVSS.n1399 DVSS 0.0148581
R10764 DVSS.n1398 DVSS 0.0148581
R10765 DVSS DVSS.n1406 0.0148581
R10766 DVSS DVSS.n1407 0.0148581
R10767 DVSS.n1420 DVSS.n1419 0.0148581
R10768 DVSS.n1422 DVSS 0.0148581
R10769 DVSS.n1421 DVSS 0.0148581
R10770 DVSS DVSS.n1432 0.0148581
R10771 DVSS DVSS.n1433 0.0148581
R10772 DVSS.n1435 DVSS 0.0148581
R10773 DVSS.n1434 DVSS 0.0148581
R10774 DVSS DVSS.n1444 0.0148581
R10775 DVSS.n1447 DVSS 0.0148581
R10776 DVSS DVSS.n1450 0.0148581
R10777 DVSS.n1452 DVSS 0.0148581
R10778 DVSS.n1451 DVSS 0.0148581
R10779 DVSS DVSS.n1459 0.0148581
R10780 DVSS DVSS.n1460 0.0148581
R10781 DVSS.n1468 DVSS 0.0148581
R10782 DVSS.n1467 DVSS 0.0148581
R10783 DVSS.n1466 DVSS 0.0148581
R10784 DVSS DVSS.n1476 0.0148581
R10785 DVSS.n1478 DVSS 0.0148581
R10786 DVSS.n1477 DVSS 0.0148581
R10787 DVSS.n1485 DVSS 0.0148581
R10788 DVSS.n1484 DVSS 0.0148581
R10789 DVSS DVSS.n1481 0.0148581
R10790 DVSS.n1482 DVSS 0.0148581
R10791 DVSS DVSS.n1493 0.0148581
R10792 DVSS DVSS.n1494 0.0148581
R10793 DVSS.n1496 DVSS 0.0148581
R10794 DVSS.n1495 DVSS 0.0148581
R10795 DVSS.n1512 DVSS.n556 0.0148581
R10796 DVSS DVSS.n1521 0.0148581
R10797 DVSS DVSS.n1522 0.0148581
R10798 DVSS.n1647 DVSS 0.0148581
R10799 DVSS.n1646 DVSS 0.0148581
R10800 DVSS.n1645 DVSS 0.0148581
R10801 DVSS.n1642 DVSS 0.0148581
R10802 DVSS.n1641 DVSS 0.0148581
R10803 DVSS.n1640 DVSS 0.0148581
R10804 DVSS DVSS.n1531 0.0148581
R10805 DVSS.n1633 DVSS 0.0148581
R10806 DVSS.n1632 DVSS 0.0148581
R10807 DVSS.n1631 DVSS 0.0148581
R10808 DVSS.n1535 DVSS 0.0148581
R10809 DVSS DVSS.n1539 0.0148581
R10810 DVSS.n1540 DVSS 0.0148581
R10811 DVSS.n1623 DVSS 0.0148581
R10812 DVSS.n1622 DVSS 0.0148581
R10813 DVSS.n1546 DVSS 0.0148581
R10814 DVSS.n1619 DVSS 0.0148581
R10815 DVSS.n1618 DVSS 0.0148581
R10816 DVSS.n1617 DVSS 0.0148581
R10817 DVSS.n1549 DVSS 0.0148581
R10818 DVSS.n1615 DVSS 0.0148581
R10819 DVSS.n1614 DVSS 0.0148581
R10820 DVSS.n1611 DVSS 0.0148581
R10821 DVSS.n1610 DVSS 0.0148581
R10822 DVSS.n1609 DVSS 0.0148581
R10823 DVSS.n1596 DVSS.n1560 0.0148581
R10824 DVSS.n1595 DVSS 0.0148581
R10825 DVSS.n1594 DVSS 0.0148581
R10826 DVSS.n1564 DVSS 0.0148581
R10827 DVSS DVSS.n1844 0.0148581
R10828 DVSS DVSS.n1845 0.0148581
R10829 DVSS.n1847 DVSS 0.0148581
R10830 DVSS.n1846 DVSS 0.0148581
R10831 DVSS.n1857 DVSS 0.0148581
R10832 DVSS DVSS.n1860 0.0148581
R10833 DVSS DVSS.n1861 0.0148581
R10834 DVSS.n1864 DVSS 0.0148581
R10835 DVSS.n1863 DVSS 0.0148581
R10836 DVSS.n1862 DVSS 0.0148581
R10837 DVSS.n1873 DVSS 0.0148581
R10838 DVSS.n1879 DVSS 0.0148581
R10839 DVSS.n1878 DVSS 0.0148581
R10840 DVSS.n462 DVSS 0.0148581
R10841 DVSS.n1888 DVSS 0.0148581
R10842 DVSS.n1887 DVSS 0.0148581
R10843 DVSS.n458 DVSS 0.0148581
R10844 DVSS.n455 DVSS 0.0148581
R10845 DVSS.n1893 DVSS 0.0148581
R10846 DVSS.n1892 DVSS 0.0148581
R10847 DVSS.n453 DVSS 0.0148581
R10848 DVSS DVSS.n1901 0.0148581
R10849 DVSS DVSS.n1902 0.0148581
R10850 DVSS.n1903 DVSS 0.0148581
R10851 DVSS.n1921 DVSS.n444 0.0148581
R10852 DVSS DVSS.n1922 0.0148581
R10853 DVSS.n1924 DVSS 0.0148581
R10854 DVSS.n1923 DVSS 0.0148581
R10855 DVSS DVSS.n2026 0.0148581
R10856 DVSS DVSS.n2027 0.0148581
R10857 DVSS.n2029 DVSS 0.0148581
R10858 DVSS.n2028 DVSS 0.0148581
R10859 DVSS.n2039 DVSS 0.0148581
R10860 DVSS DVSS.n2042 0.0148581
R10861 DVSS DVSS.n2043 0.0148581
R10862 DVSS.n2046 DVSS 0.0148581
R10863 DVSS.n2045 DVSS 0.0148581
R10864 DVSS.n2044 DVSS 0.0148581
R10865 DVSS.n2055 DVSS 0.0148581
R10866 DVSS.n2061 DVSS 0.0148581
R10867 DVSS.n2060 DVSS 0.0148581
R10868 DVSS.n390 DVSS 0.0148581
R10869 DVSS.n2070 DVSS 0.0148581
R10870 DVSS.n2069 DVSS 0.0148581
R10871 DVSS.n386 DVSS 0.0148581
R10872 DVSS.n383 DVSS 0.0148581
R10873 DVSS.n2075 DVSS 0.0148581
R10874 DVSS.n2074 DVSS 0.0148581
R10875 DVSS.n381 DVSS 0.0148581
R10876 DVSS DVSS.n2083 0.0148581
R10877 DVSS DVSS.n2084 0.0148581
R10878 DVSS.n2085 DVSS 0.0148581
R10879 DVSS.n2103 DVSS.n372 0.0148581
R10880 DVSS DVSS.n2104 0.0148581
R10881 DVSS.n2106 DVSS 0.0148581
R10882 DVSS.n2105 DVSS 0.0148581
R10883 DVSS DVSS.n2208 0.0148581
R10884 DVSS DVSS.n2209 0.0148581
R10885 DVSS.n2211 DVSS 0.0148581
R10886 DVSS.n2210 DVSS 0.0148581
R10887 DVSS.n2221 DVSS 0.0148581
R10888 DVSS DVSS.n2224 0.0148581
R10889 DVSS DVSS.n2225 0.0148581
R10890 DVSS.n2228 DVSS 0.0148581
R10891 DVSS.n2227 DVSS 0.0148581
R10892 DVSS.n2226 DVSS 0.0148581
R10893 DVSS.n2237 DVSS 0.0148581
R10894 DVSS.n2243 DVSS 0.0148581
R10895 DVSS.n2242 DVSS 0.0148581
R10896 DVSS.n318 DVSS 0.0148581
R10897 DVSS.n2252 DVSS 0.0148581
R10898 DVSS.n2251 DVSS 0.0148581
R10899 DVSS.n314 DVSS 0.0148581
R10900 DVSS.n311 DVSS 0.0148581
R10901 DVSS.n2257 DVSS 0.0148581
R10902 DVSS.n2256 DVSS 0.0148581
R10903 DVSS.n309 DVSS 0.0148581
R10904 DVSS DVSS.n2265 0.0148581
R10905 DVSS DVSS.n2266 0.0148581
R10906 DVSS.n2267 DVSS 0.0148581
R10907 DVSS.n2285 DVSS.n300 0.0148581
R10908 DVSS DVSS.n2286 0.0148581
R10909 DVSS.n2288 DVSS 0.0148581
R10910 DVSS.n2287 DVSS 0.0148581
R10911 DVSS DVSS.n2379 0.0148581
R10912 DVSS DVSS.n2380 0.0148581
R10913 DVSS.n2382 DVSS 0.0148581
R10914 DVSS.n2381 DVSS 0.0148581
R10915 DVSS.n2393 DVSS 0.0148581
R10916 DVSS DVSS.n2396 0.0148581
R10917 DVSS DVSS.n2397 0.0148581
R10918 DVSS.n2400 DVSS 0.0148581
R10919 DVSS.n2399 DVSS 0.0148581
R10920 DVSS.n2398 DVSS 0.0148581
R10921 DVSS.n2409 DVSS 0.0148581
R10922 DVSS.n2415 DVSS 0.0148581
R10923 DVSS.n2414 DVSS 0.0148581
R10924 DVSS.n117 DVSS 0.0148581
R10925 DVSS.n2427 DVSS 0.0148581
R10926 DVSS.n2426 DVSS 0.0148581
R10927 DVSS.n2423 DVSS 0.0148581
R10928 DVSS.n111 DVSS 0.0148581
R10929 DVSS.n110 DVSS 0.0148581
R10930 DVSS DVSS.n2431 0.0148581
R10931 DVSS.n2433 DVSS 0.0148581
R10932 DVSS.n2432 DVSS 0.0148581
R10933 DVSS DVSS.n2440 0.0148581
R10934 DVSS DVSS.n2441 0.0148581
R10935 DVSS.n2454 DVSS.n2453 0.0148581
R10936 DVSS.n2456 DVSS 0.0148581
R10937 DVSS.n2455 DVSS 0.0148581
R10938 DVSS DVSS.n2466 0.0148581
R10939 DVSS DVSS.n2467 0.0148581
R10940 DVSS.n2469 DVSS 0.0148581
R10941 DVSS.n2468 DVSS 0.0148581
R10942 DVSS DVSS.n2478 0.0148581
R10943 DVSS.n2481 DVSS 0.0148581
R10944 DVSS DVSS.n2484 0.0148581
R10945 DVSS.n2486 DVSS 0.0148581
R10946 DVSS.n2485 DVSS 0.0148581
R10947 DVSS DVSS.n2493 0.0148581
R10948 DVSS DVSS.n2494 0.0148581
R10949 DVSS.n2502 DVSS 0.0148581
R10950 DVSS.n2501 DVSS 0.0148581
R10951 DVSS.n2500 DVSS 0.0148581
R10952 DVSS DVSS.n2510 0.0148581
R10953 DVSS.n2512 DVSS 0.0148581
R10954 DVSS.n2511 DVSS 0.0148581
R10955 DVSS.n2519 DVSS 0.0148581
R10956 DVSS.n2518 DVSS 0.0148581
R10957 DVSS DVSS.n2515 0.0148581
R10958 DVSS.n2516 DVSS 0.0148581
R10959 DVSS DVSS.n2527 0.0148581
R10960 DVSS DVSS.n2528 0.0148581
R10961 DVSS.n2530 DVSS 0.0148581
R10962 DVSS.n2529 DVSS 0.0148581
R10963 DVSS.n2546 DVSS.n64 0.0148581
R10964 DVSS DVSS.n2555 0.0148581
R10965 DVSS DVSS.n2556 0.0148581
R10966 DVSS.n2640 DVSS 0.0148581
R10967 DVSS.n2639 DVSS 0.0148581
R10968 DVSS.n2638 DVSS 0.0148581
R10969 DVSS.n2635 DVSS 0.0148581
R10970 DVSS.n2634 DVSS 0.0148581
R10971 DVSS.n2633 DVSS 0.0148581
R10972 DVSS DVSS.n2571 0.0148581
R10973 DVSS.n2626 DVSS 0.0148581
R10974 DVSS.n2625 DVSS 0.0148581
R10975 DVSS.n2624 DVSS 0.0148581
R10976 DVSS.n2577 DVSS 0.0148581
R10977 DVSS DVSS.n2581 0.0148581
R10978 DVSS.n2582 DVSS 0.0148581
R10979 DVSS.n2616 DVSS 0.0148581
R10980 DVSS.n2615 DVSS 0.0148581
R10981 DVSS.n2592 DVSS 0.0148581
R10982 DVSS.n2612 DVSS 0.0148581
R10983 DVSS.n2611 DVSS 0.0148581
R10984 DVSS.n2610 DVSS 0.0148581
R10985 DVSS.n2595 DVSS 0.0148581
R10986 DVSS.n2608 DVSS 0.0148581
R10987 DVSS.n2607 DVSS 0.0148581
R10988 DVSS.n2604 DVSS 0.0148581
R10989 DVSS.n2603 DVSS 0.0148581
R10990 DVSS DVSS.n2787 0.0148581
R10991 DVSS.n1022 DVSS 0.0140135
R10992 DVSS.n1204 DVSS 0.0140135
R10993 DVSS.n1376 DVSS 0.0140135
R10994 DVSS.n1462 DVSS 0.0140135
R10995 DVSS.n1627 DVSS 0.0140135
R10996 DVSS.n1874 DVSS 0.0140135
R10997 DVSS.n2056 DVSS 0.0140135
R10998 DVSS.n2238 DVSS 0.0140135
R10999 DVSS.n2410 DVSS 0.0140135
R11000 DVSS.n2496 DVSS 0.0140135
R11001 DVSS.n2620 DVSS 0.0140135
R11002 DVSS.n1116 DVSS 0.0123243
R11003 DVSS.n1298 DVSS 0.0123243
R11004 DVSS DVSS.n735 0.0123243
R11005 DVSS DVSS.n1688 0.0123243
R11006 DVSS.n1786 DVSS 0.0123243
R11007 DVSS.n1968 DVSS 0.0123243
R11008 DVSS.n2150 DVSS 0.0123243
R11009 DVSS.n2332 DVSS 0.0123243
R11010 DVSS DVSS.n243 0.0123243
R11011 DVSS DVSS.n2681 0.0123243
R11012 DVSS DVSS.n2765 0.0123243
R11013 DVSS.n960 DVSS 0.0114797
R11014 DVSS.n977 DVSS 0.0114797
R11015 DVSS.n1142 DVSS 0.0114797
R11016 DVSS.n1159 DVSS 0.0114797
R11017 DVSS.n1324 DVSS 0.0114797
R11018 DVSS.n1330 DVSS 0.0114797
R11019 DVSS.n717 DVSS 0.0114797
R11020 DVSS.n707 DVSS 0.0114797
R11021 DVSS.n1741 DVSS 0.0114797
R11022 DVSS.n1731 DVSS 0.0114797
R11023 DVSS.n1812 DVSS 0.0114797
R11024 DVSS.n1829 DVSS 0.0114797
R11025 DVSS.n1994 DVSS 0.0114797
R11026 DVSS.n2011 DVSS 0.0114797
R11027 DVSS.n2176 DVSS 0.0114797
R11028 DVSS.n2193 DVSS 0.0114797
R11029 DVSS.n2358 DVSS 0.0114797
R11030 DVSS.n2364 DVSS 0.0114797
R11031 DVSS.n225 DVSS 0.0114797
R11032 DVSS.n215 DVSS 0.0114797
R11033 DVSS.n2734 DVSS 0.0114797
R11034 DVSS.n2724 DVSS 0.0114797
R11035 DVSS.n1009 DVSS 0.0114797
R11036 DVSS.n1191 DVSS 0.0114797
R11037 DVSS.n1363 DVSS 0.0114797
R11038 DVSS.n1452 DVSS 0.0114797
R11039 DVSS.n1633 DVSS 0.0114797
R11040 DVSS.n1861 DVSS 0.0114797
R11041 DVSS.n2043 DVSS 0.0114797
R11042 DVSS.n2225 DVSS 0.0114797
R11043 DVSS.n2397 DVSS 0.0114797
R11044 DVSS.n2486 DVSS 0.0114797
R11045 DVSS.n2626 DVSS 0.0114797
R11046 DVSS.n935 DVSS.n933 0.0106351
R11047 DVSS.n1058 DVSS.n1056 0.0106351
R11048 DVSS.n1240 DVSS.n1238 0.0106351
R11049 DVSS.n1408 DVSS.n594 0.0106351
R11050 DVSS.n1506 DVSS.n1504 0.0106351
R11051 DVSS.n1606 DVSS.n1605 0.0106351
R11052 DVSS.n1910 DVSS.n1908 0.0106351
R11053 DVSS.n2092 DVSS.n2090 0.0106351
R11054 DVSS.n2274 DVSS.n2272 0.0106351
R11055 DVSS.n2442 DVSS.n102 0.0106351
R11056 DVSS.n2540 DVSS.n2538 0.0106351
R11057 DVSS.n974 DVSS 0.00979054
R11058 DVSS.n1087 DVSS 0.00979054
R11059 DVSS.n1156 DVSS 0.00979054
R11060 DVSS.n1269 DVSS 0.00979054
R11061 DVSS.n1327 DVSS 0.00979054
R11062 DVSS.n755 DVSS 0.00979054
R11063 DVSS DVSS.n709 0.00979054
R11064 DVSS.n1663 DVSS 0.00979054
R11065 DVSS.n1729 DVSS 0.00979054
R11066 DVSS.n1746 DVSS 0.00979054
R11067 DVSS.n1826 DVSS 0.00979054
R11068 DVSS.n1939 DVSS 0.00979054
R11069 DVSS.n2008 DVSS 0.00979054
R11070 DVSS.n2121 DVSS 0.00979054
R11071 DVSS.n2190 DVSS 0.00979054
R11072 DVSS.n2303 DVSS 0.00979054
R11073 DVSS.n2361 DVSS 0.00979054
R11074 DVSS.n263 DVSS 0.00979054
R11075 DVSS DVSS.n217 0.00979054
R11076 DVSS.n2656 DVSS 0.00979054
R11077 DVSS.n2722 DVSS 0.00979054
R11078 DVSS.n2739 DVSS 0.00979054
R11079 DVSS.n1003 DVSS 0.00979054
R11080 DVSS.n1185 DVSS 0.00979054
R11081 DVSS.n1357 DVSS 0.00979054
R11082 DVSS.n1445 DVSS 0.00979054
R11083 DVSS.n1636 DVSS 0.00979054
R11084 DVSS.n1855 DVSS 0.00979054
R11085 DVSS.n2037 DVSS 0.00979054
R11086 DVSS.n2219 DVSS 0.00979054
R11087 DVSS.n2391 DVSS 0.00979054
R11088 DVSS.n2479 DVSS 0.00979054
R11089 DVSS.n2629 DVSS 0.00979054
R11090 DVSS.n1112 DVSS 0.00894595
R11091 DVSS.n1294 DVSS 0.00894595
R11092 DVSS DVSS.n645 0.00894595
R11093 DVSS.n1693 DVSS 0.00894595
R11094 DVSS.n1782 DVSS 0.00894595
R11095 DVSS.n1964 DVSS 0.00894595
R11096 DVSS.n2146 DVSS 0.00894595
R11097 DVSS.n2328 DVSS 0.00894595
R11098 DVSS DVSS.n153 0.00894595
R11099 DVSS.n2686 DVSS 0.00894595
R11100 DVSS.n2770 DVSS 0.00894595
R11101 DVSS DVSS.n1010 0.00725676
R11102 DVSS.n1036 DVSS 0.00725676
R11103 DVSS DVSS.n1192 0.00725676
R11104 DVSS.n1218 DVSS 0.00725676
R11105 DVSS DVSS.n1364 0.00725676
R11106 DVSS.n1393 DVSS 0.00725676
R11107 DVSS.n1460 DVSS 0.00725676
R11108 DVSS.n1478 DVSS 0.00725676
R11109 DVSS.n1535 DVSS 0.00725676
R11110 DVSS.n1546 DVSS 0.00725676
R11111 DVSS DVSS.n1862 0.00725676
R11112 DVSS.n1888 DVSS 0.00725676
R11113 DVSS DVSS.n2044 0.00725676
R11114 DVSS.n2070 DVSS 0.00725676
R11115 DVSS DVSS.n2226 0.00725676
R11116 DVSS.n2252 DVSS 0.00725676
R11117 DVSS DVSS.n2398 0.00725676
R11118 DVSS.n2427 DVSS 0.00725676
R11119 DVSS.n2494 DVSS 0.00725676
R11120 DVSS.n2512 DVSS 0.00725676
R11121 DVSS.n2577 DVSS 0.00725676
R11122 DVSS.n2592 DVSS 0.00725676
R11123 DVSS.n1113 DVSS.n1112 0.00641216
R11124 DVSS.n1295 DVSS.n1294 0.00641216
R11125 DVSS.n740 DVSS.n645 0.00641216
R11126 DVSS.n1693 DVSS.n1687 0.00641216
R11127 DVSS.n1783 DVSS.n1782 0.00641216
R11128 DVSS.n1965 DVSS.n1964 0.00641216
R11129 DVSS.n2147 DVSS.n2146 0.00641216
R11130 DVSS.n2329 DVSS.n2328 0.00641216
R11131 DVSS.n248 DVSS.n153 0.00641216
R11132 DVSS.n2686 DVSS.n2680 0.00641216
R11133 DVSS.n2770 DVSS.n2761 0.00641216
R11134 DVSS.n2762 DVSS 0.00556757
R11135 DVSS.n1004 DVSS.n1003 0.00556757
R11136 DVSS.n1041 DVSS 0.00556757
R11137 DVSS.n1186 DVSS.n1185 0.00556757
R11138 DVSS.n1223 DVSS 0.00556757
R11139 DVSS.n1358 DVSS.n1357 0.00556757
R11140 DVSS DVSS.n602 0.00556757
R11141 DVSS.n1446 DVSS.n1445 0.00556757
R11142 DVSS.n1481 DVSS 0.00556757
R11143 DVSS.n1637 DVSS.n1636 0.00556757
R11144 DVSS.n1549 DVSS 0.00556757
R11145 DVSS.n1856 DVSS.n1855 0.00556757
R11146 DVSS.n1893 DVSS 0.00556757
R11147 DVSS.n2038 DVSS.n2037 0.00556757
R11148 DVSS.n2075 DVSS 0.00556757
R11149 DVSS.n2220 DVSS.n2219 0.00556757
R11150 DVSS.n2257 DVSS 0.00556757
R11151 DVSS.n2392 DVSS.n2391 0.00556757
R11152 DVSS DVSS.n110 0.00556757
R11153 DVSS.n2480 DVSS.n2479 0.00556757
R11154 DVSS.n2515 DVSS 0.00556757
R11155 DVSS.n2630 DVSS.n2629 0.00556757
R11156 DVSS.n2595 DVSS 0.00556757
R11157 DVSS.n960 DVSS.n959 0.00387838
R11158 DVSS.n978 DVSS.n977 0.00387838
R11159 DVSS.n1142 DVSS.n1141 0.00387838
R11160 DVSS.n1160 DVSS.n1159 0.00387838
R11161 DVSS.n1324 DVSS.n1323 0.00387838
R11162 DVSS.n1331 DVSS.n1330 0.00387838
R11163 DVSS.n718 DVSS.n717 0.00387838
R11164 DVSS.n707 DVSS.n705 0.00387838
R11165 DVSS.n1741 DVSS.n1740 0.00387838
R11166 DVSS.n1732 DVSS.n1731 0.00387838
R11167 DVSS.n1812 DVSS.n1811 0.00387838
R11168 DVSS.n1830 DVSS.n1829 0.00387838
R11169 DVSS.n1994 DVSS.n1993 0.00387838
R11170 DVSS.n2012 DVSS.n2011 0.00387838
R11171 DVSS.n2176 DVSS.n2175 0.00387838
R11172 DVSS.n2194 DVSS.n2193 0.00387838
R11173 DVSS.n2358 DVSS.n2357 0.00387838
R11174 DVSS.n2365 DVSS.n2364 0.00387838
R11175 DVSS.n226 DVSS.n225 0.00387838
R11176 DVSS.n215 DVSS.n213 0.00387838
R11177 DVSS.n2734 DVSS.n2733 0.00387838
R11178 DVSS.n2725 DVSS.n2724 0.00387838
R11179 DVSS.n937 DVSS.n936 0.00387838
R11180 DVSS.n942 DVSS.n941 0.00387838
R11181 DVSS.n1060 DVSS.n1059 0.00387838
R11182 DVSS.n1065 DVSS.n1064 0.00387838
R11183 DVSS.n1242 DVSS.n1241 0.00387838
R11184 DVSS.n1247 DVSS.n1246 0.00387838
R11185 DVSS.n1415 DVSS.n1414 0.00387838
R11186 DVSS.n1416 DVSS.n590 0.00387838
R11187 DVSS.n1508 DVSS.n1507 0.00387838
R11188 DVSS.n1513 DVSS.n555 0.00387838
R11189 DVSS.n1601 DVSS.n1557 0.00387838
R11190 DVSS.n1600 DVSS.n1599 0.00387838
R11191 DVSS.n1912 DVSS.n1911 0.00387838
R11192 DVSS.n1917 DVSS.n1916 0.00387838
R11193 DVSS.n2094 DVSS.n2093 0.00387838
R11194 DVSS.n2099 DVSS.n2098 0.00387838
R11195 DVSS.n2276 DVSS.n2275 0.00387838
R11196 DVSS.n2281 DVSS.n2280 0.00387838
R11197 DVSS.n2449 DVSS.n2448 0.00387838
R11198 DVSS.n2450 DVSS.n98 0.00387838
R11199 DVSS.n2542 DVSS.n2541 0.00387838
R11200 DVSS.n2547 DVSS.n63 0.00387838
R11201 DVSS.n983 DVSS 0.00303378
R11202 DVSS.n1165 DVSS 0.00303378
R11203 DVSS.n1336 DVSS 0.00303378
R11204 DVSS DVSS.n714 0.00303378
R11205 DVSS.n1737 DVSS 0.00303378
R11206 DVSS.n1835 DVSS 0.00303378
R11207 DVSS.n2017 DVSS 0.00303378
R11208 DVSS.n2199 DVSS 0.00303378
R11209 DVSS.n2370 DVSS 0.00303378
R11210 DVSS DVSS.n222 0.00303378
R11211 DVSS.n2730 DVSS 0.00303378
R11212 DVSS.n1005 DVSS 0.00134459
R11213 DVSS.n1022 DVSS.n1020 0.00134459
R11214 DVSS.n1187 DVSS 0.00134459
R11215 DVSS.n1204 DVSS.n1202 0.00134459
R11216 DVSS.n1359 DVSS 0.00134459
R11217 DVSS.n1376 DVSS.n1374 0.00134459
R11218 DVSS.n1447 DVSS 0.00134459
R11219 DVSS.n1462 DVSS.n1461 0.00134459
R11220 DVSS DVSS.n1640 0.00134459
R11221 DVSS.n1628 DVSS.n1627 0.00134459
R11222 DVSS.n1857 DVSS 0.00134459
R11223 DVSS.n1874 DVSS.n1872 0.00134459
R11224 DVSS.n2039 DVSS 0.00134459
R11225 DVSS.n2056 DVSS.n2054 0.00134459
R11226 DVSS.n2221 DVSS 0.00134459
R11227 DVSS.n2238 DVSS.n2236 0.00134459
R11228 DVSS.n2393 DVSS 0.00134459
R11229 DVSS.n2410 DVSS.n2408 0.00134459
R11230 DVSS.n2481 DVSS 0.00134459
R11231 DVSS.n2496 DVSS.n2495 0.00134459
R11232 DVSS DVSS.n2633 0.00134459
R11233 DVSS.n2621 DVSS.n2620 0.00134459
R11234 D93v3.n6 D93v3.n5 873.303
R11235 D93v3 D93v3.n6 585
R11236 D93v3.t1 D93v3 506.99
R11237 D93v3 D93v3.t0 150.315
R11238 D93v3.n6 D93v3.t1 147.756
R11239 D93v3.n1 D93v3.t14 105.097
R11240 D93v3.n2 D93v3.t12 105.097
R11241 D93v3.n3 D93v3.t11 104.712
R11242 D93v3.n3 D93v3.t25 104.712
R11243 D93v3.n3 D93v3.t23 104.712
R11244 D93v3.n3 D93v3.t29 104.712
R11245 D93v3.n1 D93v3.t9 104.712
R11246 D93v3.n1 D93v3.t7 104.712
R11247 D93v3.n1 D93v3.t21 104.712
R11248 D93v3.n1 D93v3.t19 104.712
R11249 D93v3.n1 D93v3.t27 104.712
R11250 D93v3.n1 D93v3.t3 104.712
R11251 D93v3.n1 D93v3.t5 104.712
R11252 D93v3.n1 D93v3.t17 104.712
R11253 D93v3.n0 D93v3.t13 104.712
R11254 D93v3.n0 D93v3.t10 104.712
R11255 D93v3.n0 D93v3.t24 104.712
R11256 D93v3.n0 D93v3.t22 104.712
R11257 D93v3.n0 D93v3.t28 104.712
R11258 D93v3.n0 D93v3.t8 104.712
R11259 D93v3.n2 D93v3.t6 104.712
R11260 D93v3.n2 D93v3.t20 104.712
R11261 D93v3.n2 D93v3.t18 104.712
R11262 D93v3.n2 D93v3.t26 104.712
R11263 D93v3.n2 D93v3.t2 104.712
R11264 D93v3.n2 D93v3.t4 104.712
R11265 D93v3.n2 D93v3.t16 104.712
R11266 D93v3.n4 D93v3.t15 99.9875
R11267 D93v3 D93v3.n0 30.3224
R11268 D93v3.n3 D93v3 14.5286
R11269 D93v3.n0 D93v3 14.4208
R11270 D93v3.n0 D93v3.n2 7.0475
R11271 D93v3.n0 D93v3.n4 6.84478
R11272 D93v3.n5 D93v3 4.99562
R11273 D93v3.n3 D93v3.n1 4.838
R11274 D93v3.n4 D93v3.n3 4.72499
R11275 D93v3 D93v3.n5 2.70619
R11276 a_16261_n9984.n1 a_16261_n9984.t21 24.2469
R11277 a_16261_n9984.n15 a_16261_n9984.t10 21.6428
R11278 a_16261_n9984.n15 a_16261_n9984.t7 21.5736
R11279 a_16261_n9984.n16 a_16261_n9984.t4 21.5736
R11280 a_16261_n9984.n17 a_16261_n9984.t12 21.5736
R11281 a_16261_n9984.n18 a_16261_n9984.t6 21.5736
R11282 a_16261_n9984.n19 a_16261_n9984.t3 21.5736
R11283 a_16261_n9984.n20 a_16261_n9984.t1 21.5736
R11284 a_16261_n9984.n21 a_16261_n9984.t28 21.5736
R11285 a_16261_n9984.n22 a_16261_n9984.t9 21.5736
R11286 a_16261_n9984.n23 a_16261_n9984.t2 21.5736
R11287 a_16261_n9984.n24 a_16261_n9984.t13 21.5736
R11288 a_16261_n9984.n25 a_16261_n9984.t11 21.5736
R11289 a_16261_n9984.n26 a_16261_n9984.t29 21.5736
R11290 a_16261_n9984.n14 a_16261_n9984.t5 21.5736
R11291 a_16261_n9984.n13 a_16261_n9984.t8 21.5736
R11292 a_16261_n9984.n1 a_16261_n9984.n0 19.6822
R11293 a_16261_n9984.n3 a_16261_n9984.n2 19.6822
R11294 a_16261_n9984.n5 a_16261_n9984.n4 19.6822
R11295 a_16261_n9984.n7 a_16261_n9984.n6 19.6822
R11296 a_16261_n9984.n9 a_16261_n9984.n8 19.6822
R11297 a_16261_n9984.n11 a_16261_n9984.n10 19.6822
R11298 a_16261_n9984.n12 a_16261_n9984.t22 18.7631
R11299 a_16261_n9984.n0 a_16261_n9984.t16 3.75732
R11300 a_16261_n9984.n0 a_16261_n9984.t23 3.75732
R11301 a_16261_n9984.n2 a_16261_n9984.t14 3.75732
R11302 a_16261_n9984.n2 a_16261_n9984.t17 3.75732
R11303 a_16261_n9984.n4 a_16261_n9984.t25 3.75732
R11304 a_16261_n9984.n4 a_16261_n9984.t24 3.75732
R11305 a_16261_n9984.n6 a_16261_n9984.t19 3.75732
R11306 a_16261_n9984.n6 a_16261_n9984.t18 3.75732
R11307 a_16261_n9984.n8 a_16261_n9984.t27 3.75732
R11308 a_16261_n9984.n8 a_16261_n9984.t15 3.75732
R11309 a_16261_n9984.n10 a_16261_n9984.t20 3.75732
R11310 a_16261_n9984.n10 a_16261_n9984.t26 3.75732
R11311 a_16261_n9984.n12 a_16261_n9984.n11 3.21198
R11312 a_16261_n9984.t0 a_16261_n9984.n27 1.53882
R11313 a_16261_n9984.n13 a_16261_n9984.n12 0.943131
R11314 a_16261_n9984.n11 a_16261_n9984.n9 0.808313
R11315 a_16261_n9984.n9 a_16261_n9984.n7 0.80675
R11316 a_16261_n9984.n7 a_16261_n9984.n5 0.80675
R11317 a_16261_n9984.n5 a_16261_n9984.n3 0.80675
R11318 a_16261_n9984.n3 a_16261_n9984.n1 0.80675
R11319 a_16261_n9984.n14 a_16261_n9984.n13 0.0696489
R11320 a_16261_n9984.n27 a_16261_n9984.n14 0.0696489
R11321 a_16261_n9984.n27 a_16261_n9984.n26 0.0696489
R11322 a_16261_n9984.n26 a_16261_n9984.n25 0.0696489
R11323 a_16261_n9984.n25 a_16261_n9984.n24 0.0696489
R11324 a_16261_n9984.n24 a_16261_n9984.n23 0.0696489
R11325 a_16261_n9984.n23 a_16261_n9984.n22 0.0696489
R11326 a_16261_n9984.n22 a_16261_n9984.n21 0.0696489
R11327 a_16261_n9984.n21 a_16261_n9984.n20 0.0696489
R11328 a_16261_n9984.n20 a_16261_n9984.n19 0.0696489
R11329 a_16261_n9984.n19 a_16261_n9984.n18 0.0696489
R11330 a_16261_n9984.n18 a_16261_n9984.n17 0.0696489
R11331 a_16261_n9984.n17 a_16261_n9984.n16 0.0696489
R11332 a_16261_n9984.n16 a_16261_n9984.n15 0.0696489
R11333 a_16951_764.t5 a_16951_764.n1 553.975
R11334 a_16951_764.n6 a_16951_764.t5 553.975
R11335 a_16951_764.n5 a_16951_764.t6 275.969
R11336 a_16951_764.n3 a_16951_764.t7 275.969
R11337 a_16951_764.n4 a_16951_764.t4 275.877
R11338 a_16951_764.n9 a_16951_764.t3 15.8632
R11339 a_16951_764.n10 a_16951_764.n9 13.5228
R11340 a_16951_764.n9 a_16951_764.n8 5.588
R11341 a_16951_764.n7 a_16951_764.n6 2.79633
R11342 a_16951_764.n8 a_16951_764.n7 2.52001
R11343 a_16951_764.n3 a_16951_764.n0 2.34014
R11344 a_16951_764.n2 a_16951_764.n3 2.3327
R11345 a_16951_764.n2 a_16951_764.n4 2.23523
R11346 a_16951_764.n4 a_16951_764.n0 2.23295
R11347 a_16951_764.n5 a_16951_764.n2 2.04972
R11348 a_16951_764.n0 a_16951_764.n5 2.04764
R11349 a_16951_764.n10 a_16951_764.t2 1.84683
R11350 a_16951_764.t0 a_16951_764.n10 1.84683
R11351 a_16951_764.n8 a_16951_764.t1 1.73283
R11352 a_16951_764.n7 a_16951_764.n1 1.29633
R11353 a_16951_764.n6 a_16951_764.n0 0.585777
R11354 a_16951_764.n2 a_16951_764.n1 0.569287
R11355 VOUT.n3 VOUT.t34 21.5504
R11356 VOUT.n35 VOUT.t29 21.4815
R11357 VOUT.n3 VOUT.t18 21.4809
R11358 VOUT.n4 VOUT.t19 21.4809
R11359 VOUT.n5 VOUT.t36 21.4809
R11360 VOUT.n6 VOUT.t13 21.4809
R11361 VOUT.n7 VOUT.t20 21.4809
R11362 VOUT.n8 VOUT.t27 21.4809
R11363 VOUT.n9 VOUT.t9 21.4809
R11364 VOUT.n10 VOUT.t21 21.4809
R11365 VOUT.n11 VOUT.t22 21.4809
R11366 VOUT.n12 VOUT.t24 21.4809
R11367 VOUT.n33 VOUT.t7 21.4809
R11368 VOUT.n32 VOUT.t25 21.4809
R11369 VOUT.n31 VOUT.t2 21.4809
R11370 VOUT.n30 VOUT.t3 21.4809
R11371 VOUT.n29 VOUT.t15 21.4809
R11372 VOUT.n28 VOUT.t11 21.4809
R11373 VOUT.n27 VOUT.t17 21.4809
R11374 VOUT.n26 VOUT.t10 21.4809
R11375 VOUT.n25 VOUT.t35 21.4809
R11376 VOUT.n24 VOUT.t12 21.4809
R11377 VOUT.n23 VOUT.t28 21.4809
R11378 VOUT.n22 VOUT.t37 21.4809
R11379 VOUT.n21 VOUT.t0 21.4809
R11380 VOUT.n20 VOUT.t8 21.4809
R11381 VOUT.n19 VOUT.t16 21.4809
R11382 VOUT.n18 VOUT.t26 21.4809
R11383 VOUT.n17 VOUT.t1 21.4809
R11384 VOUT.n16 VOUT.t4 21.4809
R11385 VOUT.n15 VOUT.t23 21.4809
R11386 VOUT.n14 VOUT.t14 21.4809
R11387 VOUT.n13 VOUT.t5 21.4809
R11388 VOUT.n2 VOUT.n0 13.4669
R11389 VOUT.n2 VOUT.n1 13.3799
R11390 VOUT.n36 VOUT.n35 5.29502
R11391 VOUT.n36 VOUT.t6 4.35292
R11392 VOUT VOUT.n38 2.58592
R11393 VOUT.n37 VOUT.n36 2.49267
R11394 VOUT.n38 VOUT.n2 2.00817
R11395 VOUT.n0 VOUT.t31 1.45813
R11396 VOUT.n0 VOUT.t32 1.45813
R11397 VOUT.n1 VOUT.t30 1.45813
R11398 VOUT.n1 VOUT.t33 1.45813
R11399 VOUT.n37 VOUT 0.701375
R11400 VOUT.n13 VOUT 0.696143
R11401 VOUT.n38 VOUT.n37 0.39493
R11402 VOUT.n21 VOUT.n20 0.223778
R11403 VOUT.n17 VOUT.n16 0.205963
R11404 VOUT.n29 VOUT.n28 0.196462
R11405 VOUT.n15 VOUT.n14 0.188148
R11406 VOUT.n35 VOUT.n34 0.182804
R11407 VOUT.n14 VOUT.n13 0.15727
R11408 VOUT.n4 VOUT.n3 0.0699774
R11409 VOUT.n5 VOUT.n4 0.0699774
R11410 VOUT.n6 VOUT.n5 0.0699774
R11411 VOUT.n7 VOUT.n6 0.0699774
R11412 VOUT.n8 VOUT.n7 0.0699774
R11413 VOUT.n9 VOUT.n8 0.0699774
R11414 VOUT.n10 VOUT.n9 0.0699774
R11415 VOUT.n11 VOUT.n10 0.0699774
R11416 VOUT.n12 VOUT.n11 0.0699774
R11417 VOUT.n33 VOUT.n32 0.0699774
R11418 VOUT.n32 VOUT.n31 0.0699774
R11419 VOUT.n31 VOUT.n30 0.0699774
R11420 VOUT.n30 VOUT.n29 0.0699774
R11421 VOUT.n28 VOUT.n27 0.0699774
R11422 VOUT.n27 VOUT.n26 0.0699774
R11423 VOUT.n26 VOUT.n25 0.0699774
R11424 VOUT.n25 VOUT.n24 0.0699774
R11425 VOUT.n24 VOUT.n23 0.0699774
R11426 VOUT.n23 VOUT.n22 0.0699774
R11427 VOUT.n22 VOUT.n21 0.0699774
R11428 VOUT.n20 VOUT.n19 0.0699774
R11429 VOUT.n19 VOUT.n18 0.0699774
R11430 VOUT.n18 VOUT.n17 0.0699774
R11431 VOUT.n16 VOUT.n15 0.0699774
R11432 VOUT.n34 VOUT.n33 0.0393955
R11433 VOUT.n34 VOUT.n12 0.0310819
R11434 DVDD.n8 DVDD.n6 307.762
R11435 DVDD.n119 DVDD.n11 307.76
R11436 DVDD.n115 DVDD.n18 307.76
R11437 DVDD.n111 DVDD.n25 307.76
R11438 DVDD.n107 DVDD.n32 307.76
R11439 DVDD.n103 DVDD.n39 307.76
R11440 DVDD.n99 DVDD.n46 307.76
R11441 DVDD.n95 DVDD.n53 307.76
R11442 DVDD.n91 DVDD.n60 307.76
R11443 DVDD.n87 DVDD.n67 307.76
R11444 DVDD.n83 DVDD.n74 307.76
R11445 DVDD.n4 DVDD.n1 185
R11446 DVDD.n1 DVDD.n0 185
R11447 DVDD.n16 DVDD.n13 185
R11448 DVDD.n13 DVDD.n12 185
R11449 DVDD.n23 DVDD.n20 185
R11450 DVDD.n20 DVDD.n19 185
R11451 DVDD.n30 DVDD.n27 185
R11452 DVDD.n27 DVDD.n26 185
R11453 DVDD.n37 DVDD.n34 185
R11454 DVDD.n34 DVDD.n33 185
R11455 DVDD.n44 DVDD.n41 185
R11456 DVDD.n41 DVDD.n40 185
R11457 DVDD.n51 DVDD.n48 185
R11458 DVDD.n48 DVDD.n47 185
R11459 DVDD.n58 DVDD.n55 185
R11460 DVDD.n55 DVDD.n54 185
R11461 DVDD.n65 DVDD.n62 185
R11462 DVDD.n62 DVDD.n61 185
R11463 DVDD.n72 DVDD.n69 185
R11464 DVDD.n69 DVDD.n68 185
R11465 DVDD.n79 DVDD.n76 185
R11466 DVDD.n76 DVDD.n75 185
R11467 DVDD.n2 DVDD.t24 129.546
R11468 DVDD.n14 DVDD.t36 129.546
R11469 DVDD.n21 DVDD.t0 129.546
R11470 DVDD.n28 DVDD.t6 129.546
R11471 DVDD.n35 DVDD.t12 129.546
R11472 DVDD.n42 DVDD.t34 129.546
R11473 DVDD.n49 DVDD.t40 129.546
R11474 DVDD.n56 DVDD.t18 129.546
R11475 DVDD.n63 DVDD.t38 129.546
R11476 DVDD.n70 DVDD.t22 129.546
R11477 DVDD.n77 DVDD.t30 129.546
R11478 DVDD.n5 DVDD.n0 101.644
R11479 DVDD.n17 DVDD.n12 101.644
R11480 DVDD.n24 DVDD.n19 101.644
R11481 DVDD.n31 DVDD.n26 101.644
R11482 DVDD.n38 DVDD.n33 101.644
R11483 DVDD.n45 DVDD.n40 101.644
R11484 DVDD.n52 DVDD.n47 101.644
R11485 DVDD.n59 DVDD.n54 101.644
R11486 DVDD.n66 DVDD.n61 101.644
R11487 DVDD.n73 DVDD.n68 101.644
R11488 DVDD.n80 DVDD.n75 101.644
R11489 DVDD.n5 DVDD.n4 92.5005
R11490 DVDD.n17 DVDD.n16 92.5005
R11491 DVDD.n24 DVDD.n23 92.5005
R11492 DVDD.n31 DVDD.n30 92.5005
R11493 DVDD.n38 DVDD.n37 92.5005
R11494 DVDD.n45 DVDD.n44 92.5005
R11495 DVDD.n52 DVDD.n51 92.5005
R11496 DVDD.n59 DVDD.n58 92.5005
R11497 DVDD.n66 DVDD.n65 92.5005
R11498 DVDD.n73 DVDD.n72 92.5005
R11499 DVDD.n80 DVDD.n79 92.5005
R11500 DVDD.n3 DVDD.n2 77.057
R11501 DVDD.n15 DVDD.n14 77.057
R11502 DVDD.n22 DVDD.n21 77.057
R11503 DVDD.n29 DVDD.n28 77.057
R11504 DVDD.n36 DVDD.n35 77.057
R11505 DVDD.n43 DVDD.n42 77.057
R11506 DVDD.n50 DVDD.n49 77.057
R11507 DVDD.n57 DVDD.n56 77.057
R11508 DVDD.n64 DVDD.n63 77.057
R11509 DVDD.n71 DVDD.n70 77.057
R11510 DVDD.n78 DVDD.n77 77.057
R11511 DVDD.t24 DVDD.n1 67.8576
R11512 DVDD.t36 DVDD.n13 67.8576
R11513 DVDD.t0 DVDD.n20 67.8576
R11514 DVDD.t6 DVDD.n27 67.8576
R11515 DVDD.t12 DVDD.n34 67.8576
R11516 DVDD.t34 DVDD.n41 67.8576
R11517 DVDD.t40 DVDD.n48 67.8576
R11518 DVDD.t18 DVDD.n55 67.8576
R11519 DVDD.t38 DVDD.n62 67.8576
R11520 DVDD.t22 DVDD.n69 67.8576
R11521 DVDD.t30 DVDD.n76 67.8576
R11522 DVDD.n2 DVDD.t42 47.2949
R11523 DVDD.n14 DVDD.t28 47.2949
R11524 DVDD.n21 DVDD.t8 47.2949
R11525 DVDD.n28 DVDD.t10 47.2949
R11526 DVDD.n35 DVDD.t16 47.2949
R11527 DVDD.n42 DVDD.t20 47.2949
R11528 DVDD.n49 DVDD.t4 47.2949
R11529 DVDD.n56 DVDD.t26 47.2949
R11530 DVDD.n63 DVDD.t14 47.2949
R11531 DVDD.n70 DVDD.t2 47.2949
R11532 DVDD.n77 DVDD.t32 47.2949
R11533 DVDD.n6 DVDD.t43 32.8338
R11534 DVDD.n6 DVDD.t25 32.8338
R11535 DVDD.n11 DVDD.t29 32.8338
R11536 DVDD.n11 DVDD.t37 32.8338
R11537 DVDD.n18 DVDD.t9 32.8338
R11538 DVDD.n18 DVDD.t1 32.8338
R11539 DVDD.n25 DVDD.t11 32.8338
R11540 DVDD.n25 DVDD.t7 32.8338
R11541 DVDD.n32 DVDD.t17 32.8338
R11542 DVDD.n32 DVDD.t13 32.8338
R11543 DVDD.n39 DVDD.t21 32.8338
R11544 DVDD.n39 DVDD.t35 32.8338
R11545 DVDD.n46 DVDD.t5 32.8338
R11546 DVDD.n46 DVDD.t41 32.8338
R11547 DVDD.n53 DVDD.t27 32.8338
R11548 DVDD.n53 DVDD.t19 32.8338
R11549 DVDD.n60 DVDD.t15 32.8338
R11550 DVDD.n60 DVDD.t39 32.8338
R11551 DVDD.n67 DVDD.t3 32.8338
R11552 DVDD.n67 DVDD.t23 32.8338
R11553 DVDD.n74 DVDD.t33 32.8338
R11554 DVDD.n74 DVDD.t31 32.8338
R11555 DVDD.n3 DVDD.n0 30.8889
R11556 DVDD.n4 DVDD.n3 30.8889
R11557 DVDD.n15 DVDD.n12 30.8889
R11558 DVDD.n16 DVDD.n15 30.8889
R11559 DVDD.n22 DVDD.n19 30.8889
R11560 DVDD.n23 DVDD.n22 30.8889
R11561 DVDD.n29 DVDD.n26 30.8889
R11562 DVDD.n30 DVDD.n29 30.8889
R11563 DVDD.n36 DVDD.n33 30.8889
R11564 DVDD.n37 DVDD.n36 30.8889
R11565 DVDD.n43 DVDD.n40 30.8889
R11566 DVDD.n44 DVDD.n43 30.8889
R11567 DVDD.n50 DVDD.n47 30.8889
R11568 DVDD.n51 DVDD.n50 30.8889
R11569 DVDD.n57 DVDD.n54 30.8889
R11570 DVDD.n58 DVDD.n57 30.8889
R11571 DVDD.n64 DVDD.n61 30.8889
R11572 DVDD.n65 DVDD.n64 30.8889
R11573 DVDD.n71 DVDD.n68 30.8889
R11574 DVDD.n72 DVDD.n71 30.8889
R11575 DVDD.n78 DVDD.n75 30.8889
R11576 DVDD.n79 DVDD.n78 30.8889
R11577 DVDD.n10 DVDD.n9 22.5272
R11578 DVDD.n118 DVDD.n117 22.5272
R11579 DVDD.n114 DVDD.n113 22.5272
R11580 DVDD.n110 DVDD.n109 22.5272
R11581 DVDD.n106 DVDD.n105 22.5272
R11582 DVDD.n102 DVDD.n101 22.5272
R11583 DVDD.n98 DVDD.n97 22.5272
R11584 DVDD.n94 DVDD.n93 22.5272
R11585 DVDD.n90 DVDD.n89 22.5272
R11586 DVDD.n86 DVDD.n85 22.5272
R11587 DVDD.n82 DVDD.n81 22.5272
R11588 DVDD.n9 DVDD.n8 17.4938
R11589 DVDD.n119 DVDD.n118 17.4938
R11590 DVDD.n115 DVDD.n114 17.4938
R11591 DVDD.n111 DVDD.n110 17.4938
R11592 DVDD.n107 DVDD.n106 17.4938
R11593 DVDD.n103 DVDD.n102 17.4938
R11594 DVDD.n99 DVDD.n98 17.4938
R11595 DVDD.n95 DVDD.n94 17.4938
R11596 DVDD.n91 DVDD.n90 17.4938
R11597 DVDD.n87 DVDD.n86 17.4938
R11598 DVDD.n83 DVDD.n82 17.4938
R11599 DVDD.n84 DVDD.n83 9.3005
R11600 DVDD.n88 DVDD.n87 9.3005
R11601 DVDD.n92 DVDD.n91 9.3005
R11602 DVDD.n96 DVDD.n95 9.3005
R11603 DVDD.n100 DVDD.n99 9.3005
R11604 DVDD.n104 DVDD.n103 9.3005
R11605 DVDD.n108 DVDD.n107 9.3005
R11606 DVDD.n112 DVDD.n111 9.3005
R11607 DVDD.n116 DVDD.n115 9.3005
R11608 DVDD.n120 DVDD.n119 9.3005
R11609 DVDD.n8 DVDD.n7 9.3005
R11610 DVDD.n7 DVDD 4.44575
R11611 DVDD.n9 DVDD.n5 4.32258
R11612 DVDD.n118 DVDD.n17 4.32258
R11613 DVDD.n114 DVDD.n24 4.32258
R11614 DVDD.n110 DVDD.n31 4.32258
R11615 DVDD.n106 DVDD.n38 4.32258
R11616 DVDD.n102 DVDD.n45 4.32258
R11617 DVDD.n98 DVDD.n52 4.32258
R11618 DVDD.n94 DVDD.n59 4.32258
R11619 DVDD.n90 DVDD.n66 4.32258
R11620 DVDD.n86 DVDD.n73 4.32258
R11621 DVDD.n82 DVDD.n80 4.32258
R11622 DVDD DVDD.n120 2.4391
R11623 DVDD DVDD.n116 2.4391
R11624 DVDD DVDD.n112 2.4391
R11625 DVDD DVDD.n108 2.4391
R11626 DVDD DVDD.n104 2.4391
R11627 DVDD DVDD.n100 2.4391
R11628 DVDD DVDD.n96 2.4391
R11629 DVDD DVDD.n92 2.4391
R11630 DVDD DVDD.n88 2.4391
R11631 DVDD DVDD.n84 2.4391
R11632 DVDD.n10 DVDD 0.121114
R11633 DVDD.n117 DVDD 0.121114
R11634 DVDD.n113 DVDD 0.121114
R11635 DVDD.n109 DVDD 0.121114
R11636 DVDD.n105 DVDD 0.121114
R11637 DVDD.n101 DVDD 0.121114
R11638 DVDD.n97 DVDD 0.121114
R11639 DVDD.n93 DVDD 0.121114
R11640 DVDD.n89 DVDD 0.121114
R11641 DVDD.n85 DVDD 0.121114
R11642 DVDD.n81 DVDD 0.121114
R11643 DVDD.n7 DVDD 0.0377807
R11644 DVDD DVDD.n10 0.0377807
R11645 DVDD.n120 DVDD 0.0377807
R11646 DVDD.n117 DVDD 0.0377807
R11647 DVDD.n116 DVDD 0.0377807
R11648 DVDD.n113 DVDD 0.0377807
R11649 DVDD.n112 DVDD 0.0377807
R11650 DVDD.n109 DVDD 0.0377807
R11651 DVDD.n108 DVDD 0.0377807
R11652 DVDD.n105 DVDD 0.0377807
R11653 DVDD.n104 DVDD 0.0377807
R11654 DVDD.n101 DVDD 0.0377807
R11655 DVDD.n100 DVDD 0.0377807
R11656 DVDD.n97 DVDD 0.0377807
R11657 DVDD.n96 DVDD 0.0377807
R11658 DVDD.n93 DVDD 0.0377807
R11659 DVDD.n92 DVDD 0.0377807
R11660 DVDD.n89 DVDD 0.0377807
R11661 DVDD.n88 DVDD 0.0377807
R11662 DVDD.n85 DVDD 0.0377807
R11663 DVDD.n84 DVDD 0.0377807
R11664 DVDD.n81 DVDD 0.0377807
R11665 a_16261_n4916.n1 a_16261_n4916.t18 24.2469
R11666 a_16261_n4916.n26 a_16261_n4916.t5 21.6428
R11667 a_16261_n4916.n26 a_16261_n4916.t1 21.5736
R11668 a_16261_n4916.n25 a_16261_n4916.t12 21.5736
R11669 a_16261_n4916.n24 a_16261_n4916.t2 21.5736
R11670 a_16261_n4916.n23 a_16261_n4916.t11 21.5736
R11671 a_16261_n4916.n22 a_16261_n4916.t10 21.5736
R11672 a_16261_n4916.n21 a_16261_n4916.t9 21.5736
R11673 a_16261_n4916.n20 a_16261_n4916.t3 21.5736
R11674 a_16261_n4916.n19 a_16261_n4916.t13 21.5736
R11675 a_16261_n4916.n18 a_16261_n4916.t8 21.5736
R11676 a_16261_n4916.n17 a_16261_n4916.t4 21.5736
R11677 a_16261_n4916.n16 a_16261_n4916.t29 21.5736
R11678 a_16261_n4916.n15 a_16261_n4916.t7 21.5736
R11679 a_16261_n4916.n14 a_16261_n4916.t6 21.5736
R11680 a_16261_n4916.n13 a_16261_n4916.t28 21.5736
R11681 a_16261_n4916.n1 a_16261_n4916.n0 19.6822
R11682 a_16261_n4916.n3 a_16261_n4916.n2 19.6822
R11683 a_16261_n4916.n5 a_16261_n4916.n4 19.6822
R11684 a_16261_n4916.n7 a_16261_n4916.n6 19.6822
R11685 a_16261_n4916.n9 a_16261_n4916.n8 19.6822
R11686 a_16261_n4916.n11 a_16261_n4916.n10 19.6822
R11687 a_16261_n4916.n12 a_16261_n4916.t19 18.7631
R11688 a_16261_n4916.n0 a_16261_n4916.t25 3.75732
R11689 a_16261_n4916.n0 a_16261_n4916.t20 3.75732
R11690 a_16261_n4916.n2 a_16261_n4916.t23 3.75732
R11691 a_16261_n4916.n2 a_16261_n4916.t14 3.75732
R11692 a_16261_n4916.n4 a_16261_n4916.t22 3.75732
R11693 a_16261_n4916.n4 a_16261_n4916.t21 3.75732
R11694 a_16261_n4916.n6 a_16261_n4916.t16 3.75732
R11695 a_16261_n4916.n6 a_16261_n4916.t15 3.75732
R11696 a_16261_n4916.n8 a_16261_n4916.t27 3.75732
R11697 a_16261_n4916.n8 a_16261_n4916.t24 3.75732
R11698 a_16261_n4916.n10 a_16261_n4916.t17 3.75732
R11699 a_16261_n4916.n10 a_16261_n4916.t26 3.75732
R11700 a_16261_n4916.n12 a_16261_n4916.n11 3.21198
R11701 a_16261_n4916.t0 a_16261_n4916.n27 1.53882
R11702 a_16261_n4916.n13 a_16261_n4916.n12 0.943131
R11703 a_16261_n4916.n11 a_16261_n4916.n9 0.808313
R11704 a_16261_n4916.n9 a_16261_n4916.n7 0.80675
R11705 a_16261_n4916.n7 a_16261_n4916.n5 0.80675
R11706 a_16261_n4916.n5 a_16261_n4916.n3 0.80675
R11707 a_16261_n4916.n3 a_16261_n4916.n1 0.80675
R11708 a_16261_n4916.n14 a_16261_n4916.n13 0.0696489
R11709 a_16261_n4916.n15 a_16261_n4916.n14 0.0696489
R11710 a_16261_n4916.n16 a_16261_n4916.n15 0.0696489
R11711 a_16261_n4916.n17 a_16261_n4916.n16 0.0696489
R11712 a_16261_n4916.n18 a_16261_n4916.n17 0.0696489
R11713 a_16261_n4916.n19 a_16261_n4916.n18 0.0696489
R11714 a_16261_n4916.n20 a_16261_n4916.n19 0.0696489
R11715 a_16261_n4916.n21 a_16261_n4916.n20 0.0696489
R11716 a_16261_n4916.n22 a_16261_n4916.n21 0.0696489
R11717 a_16261_n4916.n23 a_16261_n4916.n22 0.0696489
R11718 a_16261_n4916.n24 a_16261_n4916.n23 0.0696489
R11719 a_16261_n4916.n25 a_16261_n4916.n24 0.0696489
R11720 a_16261_n4916.n27 a_16261_n4916.n25 0.0696489
R11721 a_16261_n4916.n27 a_16261_n4916.n26 0.0696489
R11722 x3.R1.n151 x3.R1.t94 492.046
R11723 x3.R1.n35 x3.R1.t24 27.6402
R11724 x3.R1.n151 x3.R1.n150 26.1161
R11725 x3.R1.n152 x3.R1.n29 22.8932
R11726 x3.R1.n14 x3.R1.t26 22.474
R11727 x3.R1.n77 x3.R1.t53 21.3897
R11728 x3.R1.n2 x3.R1.n0 20.88
R11729 x3.R1.n35 x3.R1.t36 20.7069
R11730 x3.R1.n36 x3.R1.t82 20.7069
R11731 x3.R1.n37 x3.R1.t35 20.7069
R11732 x3.R1.n45 x3.R1.t0 20.7069
R11733 x3.R1.n38 x3.R1.t31 20.7059
R11734 x3.R1.n40 x3.R1.t29 20.7059
R11735 x3.R1.n41 x3.R1.t14 20.7059
R11736 x3.R1.n34 x3.R1.t37 20.7059
R11737 x3.R1.n46 x3.R1.t46 20.7059
R11738 x3.R1.n47 x3.R1.t57 20.7059
R11739 x3.R1.n32 x3.R1.t90 20.7059
R11740 x3.R1.n51 x3.R1.t83 20.7059
R11741 x3.R1.n52 x3.R1.t11 20.7059
R11742 x3.R1.n148 x3.R1.t13 20.7059
R11743 x3.R1.n147 x3.R1.t49 20.7059
R11744 x3.R1.n146 x3.R1.t30 20.7059
R11745 x3.R1.n53 x3.R1.t2 20.7059
R11746 x3.R1.n142 x3.R1.t10 20.7059
R11747 x3.R1.n141 x3.R1.t61 20.7059
R11748 x3.R1.n140 x3.R1.t34 20.7059
R11749 x3.R1.n55 x3.R1.t28 20.7059
R11750 x3.R1.n136 x3.R1.t50 20.7059
R11751 x3.R1.n135 x3.R1.t3 20.7059
R11752 x3.R1.n134 x3.R1.t52 20.7059
R11753 x3.R1.n57 x3.R1.t85 20.7059
R11754 x3.R1.n130 x3.R1.t21 20.7059
R11755 x3.R1.n129 x3.R1.t43 20.7059
R11756 x3.R1.n128 x3.R1.t86 20.7059
R11757 x3.R1.n59 x3.R1.t41 20.7059
R11758 x3.R1.n124 x3.R1.t12 20.7059
R11759 x3.R1.n123 x3.R1.t25 20.7059
R11760 x3.R1.n122 x3.R1.t45 20.7059
R11761 x3.R1.n61 x3.R1.t5 20.7059
R11762 x3.R1.n118 x3.R1.t88 20.7059
R11763 x3.R1.n117 x3.R1.t39 20.7059
R11764 x3.R1.n116 x3.R1.t7 20.7059
R11765 x3.R1.n63 x3.R1.t81 20.7059
R11766 x3.R1.n112 x3.R1.t6 20.7059
R11767 x3.R1.n111 x3.R1.t80 20.7059
R11768 x3.R1.n110 x3.R1.t47 20.7059
R11769 x3.R1.n65 x3.R1.t89 20.7059
R11770 x3.R1.n106 x3.R1.t40 20.7059
R11771 x3.R1.n105 x3.R1.t91 20.7059
R11772 x3.R1.n104 x3.R1.t1 20.7059
R11773 x3.R1.n67 x3.R1.t23 20.7059
R11774 x3.R1.n100 x3.R1.t54 20.7059
R11775 x3.R1.n99 x3.R1.t33 20.7059
R11776 x3.R1.n98 x3.R1.t19 20.7059
R11777 x3.R1.n69 x3.R1.t87 20.7059
R11778 x3.R1.n94 x3.R1.t84 20.7059
R11779 x3.R1.n93 x3.R1.t17 20.7059
R11780 x3.R1.n92 x3.R1.t4 20.7059
R11781 x3.R1.n71 x3.R1.t32 20.7059
R11782 x3.R1.n88 x3.R1.t27 20.7059
R11783 x3.R1.n87 x3.R1.t22 20.7059
R11784 x3.R1.n86 x3.R1.t38 20.7059
R11785 x3.R1.n73 x3.R1.t51 20.7059
R11786 x3.R1.n82 x3.R1.t20 20.7059
R11787 x3.R1.n81 x3.R1.t9 20.7059
R11788 x3.R1.n80 x3.R1.t93 20.7059
R11789 x3.R1.n75 x3.R1.t44 20.7059
R11790 x3.R1.n76 x3.R1.t48 20.7059
R11791 x3.R1.n18 x3.R1.n17 19.9925
R11792 x3.R1.n20 x3.R1.n19 19.9925
R11793 x3.R1.n12 x3.R1.n11 19.9842
R11794 x3.R1.n10 x3.R1.n9 19.9842
R11795 x3.R1.n8 x3.R1.n7 19.9842
R11796 x3.R1.n6 x3.R1.n5 19.9842
R11797 x3.R1.n4 x3.R1.n3 19.9842
R11798 x3.R1.n2 x3.R1.n1 19.9842
R11799 x3.R1.n22 x3.R1.n21 19.9788
R11800 x3.R1.n24 x3.R1.n23 19.9788
R11801 x3.R1.n26 x3.R1.n25 19.9788
R11802 x3.R1.n28 x3.R1.n27 19.9788
R11803 x3.R1.n16 x3.R1.n15 19.0358
R11804 x3.R1.n13 x3.R1.t92 17.8929
R11805 x3.R1.n76 x3.R1.n75 6.93383
R11806 x3.R1.n80 x3.R1.n75 6.93383
R11807 x3.R1.n81 x3.R1.n80 6.93383
R11808 x3.R1.n82 x3.R1.n81 6.93383
R11809 x3.R1.n82 x3.R1.n73 6.93383
R11810 x3.R1.n86 x3.R1.n73 6.93383
R11811 x3.R1.n87 x3.R1.n86 6.93383
R11812 x3.R1.n88 x3.R1.n87 6.93383
R11813 x3.R1.n88 x3.R1.n71 6.93383
R11814 x3.R1.n92 x3.R1.n71 6.93383
R11815 x3.R1.n93 x3.R1.n92 6.93383
R11816 x3.R1.n94 x3.R1.n93 6.93383
R11817 x3.R1.n94 x3.R1.n69 6.93383
R11818 x3.R1.n98 x3.R1.n69 6.93383
R11819 x3.R1.n99 x3.R1.n98 6.93383
R11820 x3.R1.n100 x3.R1.n99 6.93383
R11821 x3.R1.n100 x3.R1.n67 6.93383
R11822 x3.R1.n104 x3.R1.n67 6.93383
R11823 x3.R1.n105 x3.R1.n104 6.93383
R11824 x3.R1.n106 x3.R1.n105 6.93383
R11825 x3.R1.n106 x3.R1.n65 6.93383
R11826 x3.R1.n110 x3.R1.n65 6.93383
R11827 x3.R1.n111 x3.R1.n110 6.93383
R11828 x3.R1.n112 x3.R1.n111 6.93383
R11829 x3.R1.n112 x3.R1.n63 6.93383
R11830 x3.R1.n116 x3.R1.n63 6.93383
R11831 x3.R1.n117 x3.R1.n116 6.93383
R11832 x3.R1.n118 x3.R1.n117 6.93383
R11833 x3.R1.n118 x3.R1.n61 6.93383
R11834 x3.R1.n122 x3.R1.n61 6.93383
R11835 x3.R1.n123 x3.R1.n122 6.93383
R11836 x3.R1.n124 x3.R1.n123 6.93383
R11837 x3.R1.n124 x3.R1.n59 6.93383
R11838 x3.R1.n128 x3.R1.n59 6.93383
R11839 x3.R1.n129 x3.R1.n128 6.93383
R11840 x3.R1.n130 x3.R1.n129 6.93383
R11841 x3.R1.n130 x3.R1.n57 6.93383
R11842 x3.R1.n134 x3.R1.n57 6.93383
R11843 x3.R1.n135 x3.R1.n134 6.93383
R11844 x3.R1.n136 x3.R1.n135 6.93383
R11845 x3.R1.n136 x3.R1.n55 6.93383
R11846 x3.R1.n140 x3.R1.n55 6.93383
R11847 x3.R1.n141 x3.R1.n140 6.93383
R11848 x3.R1.n142 x3.R1.n141 6.93383
R11849 x3.R1.n142 x3.R1.n53 6.93383
R11850 x3.R1.n146 x3.R1.n53 6.93383
R11851 x3.R1.n147 x3.R1.n146 6.93383
R11852 x3.R1.n148 x3.R1.n147 6.93383
R11853 x3.R1.n148 x3.R1.n52 6.93383
R11854 x3.R1.n52 x3.R1.n51 6.93383
R11855 x3.R1.n51 x3.R1.n32 6.93383
R11856 x3.R1.n47 x3.R1.n32 6.93383
R11857 x3.R1.n47 x3.R1.n46 6.93383
R11858 x3.R1.n46 x3.R1.n45 6.93383
R11859 x3.R1.n45 x3.R1.n34 6.93383
R11860 x3.R1.n41 x3.R1.n34 6.93383
R11861 x3.R1.n41 x3.R1.n40 6.93383
R11862 x3.R1.n36 x3.R1.n35 6.93383
R11863 x3.R1.n37 x3.R1.n36 6.93383
R11864 x3.R1.n38 x3.R1.n37 6.93383
R11865 x3.R1.n14 x3.R1.n13 5.42932
R11866 x3.R1.n21 x3.R1.t59 3.77447
R11867 x3.R1.n21 x3.R1.t62 3.77447
R11868 x3.R1.n23 x3.R1.t64 3.77447
R11869 x3.R1.n23 x3.R1.t58 3.77447
R11870 x3.R1.n25 x3.R1.t65 3.77447
R11871 x3.R1.n25 x3.R1.t42 3.77447
R11872 x3.R1.n27 x3.R1.t63 3.77447
R11873 x3.R1.n27 x3.R1.t60 3.77447
R11874 x3.R1.n11 x3.R1.t75 3.75732
R11875 x3.R1.n11 x3.R1.t73 3.75732
R11876 x3.R1.n9 x3.R1.t69 3.75732
R11877 x3.R1.n9 x3.R1.t68 3.75732
R11878 x3.R1.n7 x3.R1.t76 3.75732
R11879 x3.R1.n7 x3.R1.t66 3.75732
R11880 x3.R1.n5 x3.R1.t70 3.75732
R11881 x3.R1.n5 x3.R1.t77 3.75732
R11882 x3.R1.n3 x3.R1.t67 3.75732
R11883 x3.R1.n3 x3.R1.t71 3.75732
R11884 x3.R1.n1 x3.R1.t78 3.75732
R11885 x3.R1.n1 x3.R1.t79 3.75732
R11886 x3.R1.n0 x3.R1.t74 3.75732
R11887 x3.R1.n0 x3.R1.t72 3.75732
R11888 x3.R1.n17 x3.R1.t16 3.55534
R11889 x3.R1.n17 x3.R1.t15 3.55534
R11890 x3.R1.n19 x3.R1.t18 3.55534
R11891 x3.R1.n19 x3.R1.t8 3.55534
R11892 x3.R1.n15 x3.R1.t55 3.39475
R11893 x3.R1.n15 x3.R1.t56 3.39475
R11894 x3.R1.n22 x3.R1.n20 1.55606
R11895 x3.R1.n18 x3.R1.n16 1.55606
R11896 x3.R1.n16 x3.R1.n14 1.55606
R11897 x3.R1.n28 x3.R1.n26 0.898069
R11898 x3.R1.n24 x3.R1.n22 0.898069
R11899 x3.R1.n20 x3.R1.n18 0.896333
R11900 x3.R1.n4 x3.R1.n2 0.896333
R11901 x3.R1.n6 x3.R1.n4 0.896333
R11902 x3.R1.n8 x3.R1.n6 0.896333
R11903 x3.R1.n12 x3.R1.n10 0.896333
R11904 x3.R1.n26 x3.R1.n24 0.894597
R11905 x3.R1.n10 x3.R1.n8 0.894597
R11906 x3.R1.n29 x3.R1.n28 0.807609
R11907 x3.R1.n42 x3.R1.n41 0.7755
R11908 x3.R1.n43 x3.R1.n34 0.7755
R11909 x3.R1.n46 x3.R1.n33 0.7755
R11910 x3.R1.n48 x3.R1.n47 0.7755
R11911 x3.R1.n49 x3.R1.n32 0.7755
R11912 x3.R1.n51 x3.R1.n50 0.7755
R11913 x3.R1.n52 x3.R1.n30 0.7755
R11914 x3.R1.n149 x3.R1.n148 0.7755
R11915 x3.R1.n147 x3.R1.n31 0.7755
R11916 x3.R1.n146 x3.R1.n145 0.7755
R11917 x3.R1.n144 x3.R1.n53 0.7755
R11918 x3.R1.n143 x3.R1.n142 0.7755
R11919 x3.R1.n141 x3.R1.n54 0.7755
R11920 x3.R1.n140 x3.R1.n139 0.7755
R11921 x3.R1.n138 x3.R1.n55 0.7755
R11922 x3.R1.n137 x3.R1.n136 0.7755
R11923 x3.R1.n135 x3.R1.n56 0.7755
R11924 x3.R1.n134 x3.R1.n133 0.7755
R11925 x3.R1.n132 x3.R1.n57 0.7755
R11926 x3.R1.n131 x3.R1.n130 0.7755
R11927 x3.R1.n129 x3.R1.n58 0.7755
R11928 x3.R1.n128 x3.R1.n127 0.7755
R11929 x3.R1.n126 x3.R1.n59 0.7755
R11930 x3.R1.n125 x3.R1.n124 0.7755
R11931 x3.R1.n123 x3.R1.n60 0.7755
R11932 x3.R1.n122 x3.R1.n121 0.7755
R11933 x3.R1.n120 x3.R1.n61 0.7755
R11934 x3.R1.n119 x3.R1.n118 0.7755
R11935 x3.R1.n117 x3.R1.n62 0.7755
R11936 x3.R1.n116 x3.R1.n115 0.7755
R11937 x3.R1.n114 x3.R1.n63 0.7755
R11938 x3.R1.n113 x3.R1.n112 0.7755
R11939 x3.R1.n111 x3.R1.n64 0.7755
R11940 x3.R1.n110 x3.R1.n109 0.7755
R11941 x3.R1.n108 x3.R1.n65 0.7755
R11942 x3.R1.n107 x3.R1.n106 0.7755
R11943 x3.R1.n105 x3.R1.n66 0.7755
R11944 x3.R1.n104 x3.R1.n103 0.7755
R11945 x3.R1.n102 x3.R1.n67 0.7755
R11946 x3.R1.n101 x3.R1.n100 0.7755
R11947 x3.R1.n99 x3.R1.n68 0.7755
R11948 x3.R1.n98 x3.R1.n97 0.7755
R11949 x3.R1.n96 x3.R1.n69 0.7755
R11950 x3.R1.n95 x3.R1.n94 0.7755
R11951 x3.R1.n93 x3.R1.n70 0.7755
R11952 x3.R1.n92 x3.R1.n91 0.7755
R11953 x3.R1.n90 x3.R1.n71 0.7755
R11954 x3.R1.n89 x3.R1.n88 0.7755
R11955 x3.R1.n87 x3.R1.n72 0.7755
R11956 x3.R1.n86 x3.R1.n85 0.7755
R11957 x3.R1.n84 x3.R1.n73 0.7755
R11958 x3.R1.n83 x3.R1.n82 0.7755
R11959 x3.R1.n81 x3.R1.n74 0.7755
R11960 x3.R1.n80 x3.R1.n79 0.7755
R11961 x3.R1.n78 x3.R1.n75 0.7755
R11962 x3.R1.n45 x3.R1.n44 0.7755
R11963 x3.R1.n39 x3.R1.n38 0.684283
R11964 x3.R1.n29 x3.R1.n12 0.672192
R11965 x3.R1.n40 x3.R1.n39 0.629383
R11966 x3.R1.n77 x3.R1.n76 0.629383
R11967 x3.R1.n13 x3.R1 0.558313
R11968 x3.R1.n42 x3.R1.n39 0.145085
R11969 x3.R1.n78 x3.R1.n77 0.145085
R11970 x3.R1.n43 x3.R1.n42 0.0682083
R11971 x3.R1.n44 x3.R1.n43 0.0682083
R11972 x3.R1.n44 x3.R1.n33 0.0682083
R11973 x3.R1.n48 x3.R1.n33 0.0682083
R11974 x3.R1.n49 x3.R1.n48 0.0682083
R11975 x3.R1.n50 x3.R1.n49 0.0682083
R11976 x3.R1.n50 x3.R1.n30 0.0682083
R11977 x3.R1.n149 x3.R1.n31 0.0682083
R11978 x3.R1.n145 x3.R1.n31 0.0682083
R11979 x3.R1.n145 x3.R1.n144 0.0682083
R11980 x3.R1.n144 x3.R1.n143 0.0682083
R11981 x3.R1.n143 x3.R1.n54 0.0682083
R11982 x3.R1.n139 x3.R1.n54 0.0682083
R11983 x3.R1.n139 x3.R1.n138 0.0682083
R11984 x3.R1.n138 x3.R1.n137 0.0682083
R11985 x3.R1.n137 x3.R1.n56 0.0682083
R11986 x3.R1.n133 x3.R1.n56 0.0682083
R11987 x3.R1.n133 x3.R1.n132 0.0682083
R11988 x3.R1.n132 x3.R1.n131 0.0682083
R11989 x3.R1.n131 x3.R1.n58 0.0682083
R11990 x3.R1.n127 x3.R1.n58 0.0682083
R11991 x3.R1.n127 x3.R1.n126 0.0682083
R11992 x3.R1.n126 x3.R1.n125 0.0682083
R11993 x3.R1.n125 x3.R1.n60 0.0682083
R11994 x3.R1.n121 x3.R1.n60 0.0682083
R11995 x3.R1.n121 x3.R1.n120 0.0682083
R11996 x3.R1.n120 x3.R1.n119 0.0682083
R11997 x3.R1.n119 x3.R1.n62 0.0682083
R11998 x3.R1.n115 x3.R1.n62 0.0682083
R11999 x3.R1.n115 x3.R1.n114 0.0682083
R12000 x3.R1.n114 x3.R1.n113 0.0682083
R12001 x3.R1.n113 x3.R1.n64 0.0682083
R12002 x3.R1.n109 x3.R1.n64 0.0682083
R12003 x3.R1.n109 x3.R1.n108 0.0682083
R12004 x3.R1.n108 x3.R1.n107 0.0682083
R12005 x3.R1.n107 x3.R1.n66 0.0682083
R12006 x3.R1.n103 x3.R1.n66 0.0682083
R12007 x3.R1.n103 x3.R1.n102 0.0682083
R12008 x3.R1.n102 x3.R1.n101 0.0682083
R12009 x3.R1.n101 x3.R1.n68 0.0682083
R12010 x3.R1.n97 x3.R1.n68 0.0682083
R12011 x3.R1.n97 x3.R1.n96 0.0682083
R12012 x3.R1.n96 x3.R1.n95 0.0682083
R12013 x3.R1.n95 x3.R1.n70 0.0682083
R12014 x3.R1.n91 x3.R1.n70 0.0682083
R12015 x3.R1.n91 x3.R1.n90 0.0682083
R12016 x3.R1.n90 x3.R1.n89 0.0682083
R12017 x3.R1.n89 x3.R1.n72 0.0682083
R12018 x3.R1.n85 x3.R1.n72 0.0682083
R12019 x3.R1.n85 x3.R1.n84 0.0682083
R12020 x3.R1.n84 x3.R1.n83 0.0682083
R12021 x3.R1.n83 x3.R1.n74 0.0682083
R12022 x3.R1.n79 x3.R1.n74 0.0682083
R12023 x3.R1.n79 x3.R1.n78 0.0682083
R12024 x3.R1 x3.R1.n152 0.063
R12025 x3.R1.n150 x3.R1.n30 0.0560556
R12026 x3.R1.n150 x3.R1.n149 0.0126528
R12027 x3.R1.n152 x3.R1.n151 0.00154167
R12028 x5.V2.n151 x5.V2.t94 491.704
R12029 x5.V2.n152 x5.V2.n29 37.6227
R12030 x5.V2.n151 x5.V2.n150 27.7136
R12031 x5.V2.n53 x5.V2.t55 27.6402
R12032 x5.V2.n22 x5.V2.t34 22.474
R12033 x5.V2.n127 x5.V2.t63 21.3897
R12034 x5.V2.n2 x5.V2.n0 20.88
R12035 x5.V2.n53 x5.V2.t43 20.7069
R12036 x5.V2.n54 x5.V2.t53 20.7069
R12037 x5.V2.n55 x5.V2.t87 20.7069
R12038 x5.V2.n120 x5.V2.t0 20.7069
R12039 x5.V2.n56 x5.V2.t88 20.7059
R12040 x5.V2.n52 x5.V2.t12 20.7059
R12041 x5.V2.n59 x5.V2.t51 20.7059
R12042 x5.V2.n60 x5.V2.t74 20.7059
R12043 x5.V2.n61 x5.V2.t2 20.7059
R12044 x5.V2.n50 x5.V2.t66 20.7059
R12045 x5.V2.n65 x5.V2.t48 20.7059
R12046 x5.V2.n66 x5.V2.t86 20.7059
R12047 x5.V2.n67 x5.V2.t4 20.7059
R12048 x5.V2.n48 x5.V2.t14 20.7059
R12049 x5.V2.n71 x5.V2.t79 20.7059
R12050 x5.V2.n72 x5.V2.t50 20.7059
R12051 x5.V2.n73 x5.V2.t46 20.7059
R12052 x5.V2.n46 x5.V2.t93 20.7059
R12053 x5.V2.n77 x5.V2.t76 20.7059
R12054 x5.V2.n78 x5.V2.t38 20.7059
R12055 x5.V2.n79 x5.V2.t42 20.7059
R12056 x5.V2.n44 x5.V2.t20 20.7059
R12057 x5.V2.n83 x5.V2.t49 20.7059
R12058 x5.V2.n84 x5.V2.t81 20.7059
R12059 x5.V2.n85 x5.V2.t89 20.7059
R12060 x5.V2.n42 x5.V2.t7 20.7059
R12061 x5.V2.n89 x5.V2.t44 20.7059
R12062 x5.V2.n90 x5.V2.t30 20.7059
R12063 x5.V2.n91 x5.V2.t54 20.7059
R12064 x5.V2.n40 x5.V2.t31 20.7059
R12065 x5.V2.n95 x5.V2.t90 20.7059
R12066 x5.V2.n96 x5.V2.t19 20.7059
R12067 x5.V2.n97 x5.V2.t67 20.7059
R12068 x5.V2.n38 x5.V2.t39 20.7059
R12069 x5.V2.n101 x5.V2.t65 20.7059
R12070 x5.V2.n102 x5.V2.t37 20.7059
R12071 x5.V2.n103 x5.V2.t69 20.7059
R12072 x5.V2.n36 x5.V2.t35 20.7059
R12073 x5.V2.n107 x5.V2.t64 20.7059
R12074 x5.V2.n108 x5.V2.t3 20.7059
R12075 x5.V2.n109 x5.V2.t27 20.7059
R12076 x5.V2.n34 x5.V2.t33 20.7059
R12077 x5.V2.n113 x5.V2.t1 20.7059
R12078 x5.V2.n114 x5.V2.t28 20.7059
R12079 x5.V2.n115 x5.V2.t45 20.7059
R12080 x5.V2.n32 x5.V2.t32 20.7059
R12081 x5.V2.n119 x5.V2.t68 20.7059
R12082 x5.V2.n148 x5.V2.t80 20.7059
R12083 x5.V2.n147 x5.V2.t72 20.7059
R12084 x5.V2.n146 x5.V2.t70 20.7059
R12085 x5.V2.n121 x5.V2.t71 20.7059
R12086 x5.V2.n142 x5.V2.t73 20.7059
R12087 x5.V2.n141 x5.V2.t15 20.7059
R12088 x5.V2.n140 x5.V2.t11 20.7059
R12089 x5.V2.n123 x5.V2.t56 20.7059
R12090 x5.V2.n136 x5.V2.t85 20.7059
R12091 x5.V2.n135 x5.V2.t52 20.7059
R12092 x5.V2.n134 x5.V2.t29 20.7059
R12093 x5.V2.n125 x5.V2.t57 20.7059
R12094 x5.V2.n130 x5.V2.t13 20.7059
R12095 x5.V2.n129 x5.V2.t6 20.7059
R12096 x5.V2.n128 x5.V2.t22 20.7059
R12097 x5.V2.n26 x5.V2.n25 19.9925
R12098 x5.V2.n28 x5.V2.n27 19.9925
R12099 x5.V2.n12 x5.V2.n11 19.9842
R12100 x5.V2.n10 x5.V2.n9 19.9842
R12101 x5.V2.n8 x5.V2.n7 19.9842
R12102 x5.V2.n6 x5.V2.n5 19.9842
R12103 x5.V2.n4 x5.V2.n3 19.9842
R12104 x5.V2.n2 x5.V2.n1 19.9842
R12105 x5.V2.n20 x5.V2.n19 19.9788
R12106 x5.V2.n18 x5.V2.n17 19.9788
R12107 x5.V2.n16 x5.V2.n15 19.9788
R12108 x5.V2.n14 x5.V2.n13 19.9788
R12109 x5.V2.n24 x5.V2.n23 19.0358
R12110 x5.V2.n21 x5.V2.t92 17.8929
R12111 x5.V2.n129 x5.V2.n128 6.93383
R12112 x5.V2.n130 x5.V2.n129 6.93383
R12113 x5.V2.n130 x5.V2.n125 6.93383
R12114 x5.V2.n134 x5.V2.n125 6.93383
R12115 x5.V2.n135 x5.V2.n134 6.93383
R12116 x5.V2.n136 x5.V2.n135 6.93383
R12117 x5.V2.n136 x5.V2.n123 6.93383
R12118 x5.V2.n140 x5.V2.n123 6.93383
R12119 x5.V2.n141 x5.V2.n140 6.93383
R12120 x5.V2.n142 x5.V2.n141 6.93383
R12121 x5.V2.n142 x5.V2.n121 6.93383
R12122 x5.V2.n146 x5.V2.n121 6.93383
R12123 x5.V2.n147 x5.V2.n146 6.93383
R12124 x5.V2.n148 x5.V2.n147 6.93383
R12125 x5.V2.n148 x5.V2.n120 6.93383
R12126 x5.V2.n120 x5.V2.n119 6.93383
R12127 x5.V2.n119 x5.V2.n32 6.93383
R12128 x5.V2.n115 x5.V2.n32 6.93383
R12129 x5.V2.n115 x5.V2.n114 6.93383
R12130 x5.V2.n114 x5.V2.n113 6.93383
R12131 x5.V2.n113 x5.V2.n34 6.93383
R12132 x5.V2.n109 x5.V2.n34 6.93383
R12133 x5.V2.n109 x5.V2.n108 6.93383
R12134 x5.V2.n108 x5.V2.n107 6.93383
R12135 x5.V2.n107 x5.V2.n36 6.93383
R12136 x5.V2.n103 x5.V2.n36 6.93383
R12137 x5.V2.n103 x5.V2.n102 6.93383
R12138 x5.V2.n102 x5.V2.n101 6.93383
R12139 x5.V2.n101 x5.V2.n38 6.93383
R12140 x5.V2.n97 x5.V2.n38 6.93383
R12141 x5.V2.n97 x5.V2.n96 6.93383
R12142 x5.V2.n96 x5.V2.n95 6.93383
R12143 x5.V2.n95 x5.V2.n40 6.93383
R12144 x5.V2.n91 x5.V2.n40 6.93383
R12145 x5.V2.n91 x5.V2.n90 6.93383
R12146 x5.V2.n90 x5.V2.n89 6.93383
R12147 x5.V2.n89 x5.V2.n42 6.93383
R12148 x5.V2.n85 x5.V2.n42 6.93383
R12149 x5.V2.n85 x5.V2.n84 6.93383
R12150 x5.V2.n84 x5.V2.n83 6.93383
R12151 x5.V2.n83 x5.V2.n44 6.93383
R12152 x5.V2.n79 x5.V2.n44 6.93383
R12153 x5.V2.n79 x5.V2.n78 6.93383
R12154 x5.V2.n78 x5.V2.n77 6.93383
R12155 x5.V2.n77 x5.V2.n46 6.93383
R12156 x5.V2.n73 x5.V2.n46 6.93383
R12157 x5.V2.n73 x5.V2.n72 6.93383
R12158 x5.V2.n72 x5.V2.n71 6.93383
R12159 x5.V2.n71 x5.V2.n48 6.93383
R12160 x5.V2.n67 x5.V2.n48 6.93383
R12161 x5.V2.n67 x5.V2.n66 6.93383
R12162 x5.V2.n66 x5.V2.n65 6.93383
R12163 x5.V2.n65 x5.V2.n50 6.93383
R12164 x5.V2.n61 x5.V2.n50 6.93383
R12165 x5.V2.n61 x5.V2.n60 6.93383
R12166 x5.V2.n60 x5.V2.n59 6.93383
R12167 x5.V2.n59 x5.V2.n52 6.93383
R12168 x5.V2.n54 x5.V2.n53 6.93383
R12169 x5.V2.n55 x5.V2.n54 6.93383
R12170 x5.V2.n56 x5.V2.n55 6.93383
R12171 x5.V2.n22 x5.V2.n21 5.42932
R12172 x5.V2.n19 x5.V2.t41 3.77447
R12173 x5.V2.n19 x5.V2.t26 3.77447
R12174 x5.V2.n17 x5.V2.t59 3.77447
R12175 x5.V2.n17 x5.V2.t17 3.77447
R12176 x5.V2.n15 x5.V2.t18 3.77447
R12177 x5.V2.n15 x5.V2.t60 3.77447
R12178 x5.V2.n13 x5.V2.t58 3.77447
R12179 x5.V2.n13 x5.V2.t16 3.77447
R12180 x5.V2.n11 x5.V2.t62 3.75732
R12181 x5.V2.n11 x5.V2.t82 3.75732
R12182 x5.V2.n9 x5.V2.t10 3.75732
R12183 x5.V2.n9 x5.V2.t21 3.75732
R12184 x5.V2.n7 x5.V2.t61 3.75732
R12185 x5.V2.n7 x5.V2.t5 3.75732
R12186 x5.V2.n5 x5.V2.t9 3.75732
R12187 x5.V2.n5 x5.V2.t8 3.75732
R12188 x5.V2.n3 x5.V2.t47 3.75732
R12189 x5.V2.n3 x5.V2.t75 3.75732
R12190 x5.V2.n1 x5.V2.t83 3.75732
R12191 x5.V2.n1 x5.V2.t84 3.75732
R12192 x5.V2.n0 x5.V2.t77 3.75732
R12193 x5.V2.n0 x5.V2.t78 3.75732
R12194 x5.V2.n25 x5.V2.t23 3.55534
R12195 x5.V2.n25 x5.V2.t25 3.55534
R12196 x5.V2.n27 x5.V2.t24 3.55534
R12197 x5.V2.n27 x5.V2.t36 3.55534
R12198 x5.V2.n23 x5.V2.t91 3.39475
R12199 x5.V2.n23 x5.V2.t40 3.39475
R12200 x5.V2.n26 x5.V2.n24 1.55606
R12201 x5.V2.n24 x5.V2.n22 1.55606
R12202 x5.V2.n14 x5.V2.n12 1.55606
R12203 x5.V2.n16 x5.V2.n14 0.898069
R12204 x5.V2.n20 x5.V2.n18 0.898069
R12205 x5.V2.n28 x5.V2.n26 0.896333
R12206 x5.V2.n4 x5.V2.n2 0.896333
R12207 x5.V2.n6 x5.V2.n4 0.896333
R12208 x5.V2.n8 x5.V2.n6 0.896333
R12209 x5.V2.n12 x5.V2.n10 0.896333
R12210 x5.V2.n10 x5.V2.n8 0.894597
R12211 x5.V2.n18 x5.V2.n16 0.894597
R12212 x5.V2.n29 x5.V2.n28 0.808139
R12213 x5.V2.n59 x5.V2.n58 0.7755
R12214 x5.V2.n60 x5.V2.n51 0.7755
R12215 x5.V2.n62 x5.V2.n61 0.7755
R12216 x5.V2.n63 x5.V2.n50 0.7755
R12217 x5.V2.n65 x5.V2.n64 0.7755
R12218 x5.V2.n66 x5.V2.n49 0.7755
R12219 x5.V2.n68 x5.V2.n67 0.7755
R12220 x5.V2.n69 x5.V2.n48 0.7755
R12221 x5.V2.n71 x5.V2.n70 0.7755
R12222 x5.V2.n72 x5.V2.n47 0.7755
R12223 x5.V2.n74 x5.V2.n73 0.7755
R12224 x5.V2.n75 x5.V2.n46 0.7755
R12225 x5.V2.n77 x5.V2.n76 0.7755
R12226 x5.V2.n78 x5.V2.n45 0.7755
R12227 x5.V2.n80 x5.V2.n79 0.7755
R12228 x5.V2.n81 x5.V2.n44 0.7755
R12229 x5.V2.n83 x5.V2.n82 0.7755
R12230 x5.V2.n84 x5.V2.n43 0.7755
R12231 x5.V2.n86 x5.V2.n85 0.7755
R12232 x5.V2.n87 x5.V2.n42 0.7755
R12233 x5.V2.n89 x5.V2.n88 0.7755
R12234 x5.V2.n90 x5.V2.n41 0.7755
R12235 x5.V2.n92 x5.V2.n91 0.7755
R12236 x5.V2.n93 x5.V2.n40 0.7755
R12237 x5.V2.n95 x5.V2.n94 0.7755
R12238 x5.V2.n96 x5.V2.n39 0.7755
R12239 x5.V2.n98 x5.V2.n97 0.7755
R12240 x5.V2.n99 x5.V2.n38 0.7755
R12241 x5.V2.n101 x5.V2.n100 0.7755
R12242 x5.V2.n102 x5.V2.n37 0.7755
R12243 x5.V2.n104 x5.V2.n103 0.7755
R12244 x5.V2.n105 x5.V2.n36 0.7755
R12245 x5.V2.n107 x5.V2.n106 0.7755
R12246 x5.V2.n108 x5.V2.n35 0.7755
R12247 x5.V2.n110 x5.V2.n109 0.7755
R12248 x5.V2.n111 x5.V2.n34 0.7755
R12249 x5.V2.n113 x5.V2.n112 0.7755
R12250 x5.V2.n114 x5.V2.n33 0.7755
R12251 x5.V2.n116 x5.V2.n115 0.7755
R12252 x5.V2.n117 x5.V2.n32 0.7755
R12253 x5.V2.n119 x5.V2.n118 0.7755
R12254 x5.V2.n149 x5.V2.n148 0.7755
R12255 x5.V2.n147 x5.V2.n31 0.7755
R12256 x5.V2.n146 x5.V2.n145 0.7755
R12257 x5.V2.n144 x5.V2.n121 0.7755
R12258 x5.V2.n143 x5.V2.n142 0.7755
R12259 x5.V2.n141 x5.V2.n122 0.7755
R12260 x5.V2.n140 x5.V2.n139 0.7755
R12261 x5.V2.n138 x5.V2.n123 0.7755
R12262 x5.V2.n137 x5.V2.n136 0.7755
R12263 x5.V2.n135 x5.V2.n124 0.7755
R12264 x5.V2.n134 x5.V2.n133 0.7755
R12265 x5.V2.n132 x5.V2.n125 0.7755
R12266 x5.V2.n131 x5.V2.n130 0.7755
R12267 x5.V2.n129 x5.V2.n126 0.7755
R12268 x5.V2.n120 x5.V2.n30 0.7755
R12269 x5.V2.n29 x5.V2.n20 0.717167
R12270 x5.V2.n57 x5.V2.n56 0.684283
R12271 x5.V2.n57 x5.V2.n52 0.629383
R12272 x5.V2.n128 x5.V2.n127 0.629383
R12273 x5.V2.n21 x5.V2 0.558313
R12274 x5.V2.n152 x5.V2.n151 0.340083
R12275 x5.V2.n58 x5.V2.n57 0.145085
R12276 x5.V2.n127 x5.V2.n126 0.145085
R12277 x5.V2.n58 x5.V2.n51 0.0682083
R12278 x5.V2.n62 x5.V2.n51 0.0682083
R12279 x5.V2.n63 x5.V2.n62 0.0682083
R12280 x5.V2.n64 x5.V2.n63 0.0682083
R12281 x5.V2.n64 x5.V2.n49 0.0682083
R12282 x5.V2.n68 x5.V2.n49 0.0682083
R12283 x5.V2.n69 x5.V2.n68 0.0682083
R12284 x5.V2.n70 x5.V2.n69 0.0682083
R12285 x5.V2.n70 x5.V2.n47 0.0682083
R12286 x5.V2.n74 x5.V2.n47 0.0682083
R12287 x5.V2.n75 x5.V2.n74 0.0682083
R12288 x5.V2.n76 x5.V2.n75 0.0682083
R12289 x5.V2.n76 x5.V2.n45 0.0682083
R12290 x5.V2.n80 x5.V2.n45 0.0682083
R12291 x5.V2.n81 x5.V2.n80 0.0682083
R12292 x5.V2.n82 x5.V2.n81 0.0682083
R12293 x5.V2.n82 x5.V2.n43 0.0682083
R12294 x5.V2.n86 x5.V2.n43 0.0682083
R12295 x5.V2.n87 x5.V2.n86 0.0682083
R12296 x5.V2.n88 x5.V2.n87 0.0682083
R12297 x5.V2.n88 x5.V2.n41 0.0682083
R12298 x5.V2.n92 x5.V2.n41 0.0682083
R12299 x5.V2.n93 x5.V2.n92 0.0682083
R12300 x5.V2.n94 x5.V2.n93 0.0682083
R12301 x5.V2.n94 x5.V2.n39 0.0682083
R12302 x5.V2.n98 x5.V2.n39 0.0682083
R12303 x5.V2.n99 x5.V2.n98 0.0682083
R12304 x5.V2.n100 x5.V2.n99 0.0682083
R12305 x5.V2.n100 x5.V2.n37 0.0682083
R12306 x5.V2.n104 x5.V2.n37 0.0682083
R12307 x5.V2.n105 x5.V2.n104 0.0682083
R12308 x5.V2.n106 x5.V2.n105 0.0682083
R12309 x5.V2.n106 x5.V2.n35 0.0682083
R12310 x5.V2.n110 x5.V2.n35 0.0682083
R12311 x5.V2.n111 x5.V2.n110 0.0682083
R12312 x5.V2.n112 x5.V2.n111 0.0682083
R12313 x5.V2.n112 x5.V2.n33 0.0682083
R12314 x5.V2.n116 x5.V2.n33 0.0682083
R12315 x5.V2.n117 x5.V2.n116 0.0682083
R12316 x5.V2.n118 x5.V2.n117 0.0682083
R12317 x5.V2.n118 x5.V2.n30 0.0682083
R12318 x5.V2.n149 x5.V2.n31 0.0682083
R12319 x5.V2.n145 x5.V2.n31 0.0682083
R12320 x5.V2.n145 x5.V2.n144 0.0682083
R12321 x5.V2.n144 x5.V2.n143 0.0682083
R12322 x5.V2.n143 x5.V2.n122 0.0682083
R12323 x5.V2.n139 x5.V2.n122 0.0682083
R12324 x5.V2.n139 x5.V2.n138 0.0682083
R12325 x5.V2.n138 x5.V2.n137 0.0682083
R12326 x5.V2.n137 x5.V2.n124 0.0682083
R12327 x5.V2.n133 x5.V2.n124 0.0682083
R12328 x5.V2.n133 x5.V2.n132 0.0682083
R12329 x5.V2.n132 x5.V2.n131 0.0682083
R12330 x5.V2.n131 x5.V2.n126 0.0682083
R12331 x5.V2 x5.V2.n152 0.0650833
R12332 x5.V2.n150 x5.V2.n149 0.0514259
R12333 x5.V2.n150 x5.V2.n30 0.0172824
R12334 x4.V2.n150 x4.V2.t94 491.704
R12335 x4.V2.n27 x4.V2.t59 22.474
R12336 x4.V2.n30 x4.V2.t64 21.4824
R12337 x4.V2.n2 x4.V2.n0 20.88
R12338 x4.V2.n62 x4.V2.t89 20.7986
R12339 x4.V2.n58 x4.V2.t13 20.7986
R12340 x4.V2.n57 x4.V2.t52 20.7986
R12341 x4.V2.n66 x4.V2.t75 20.7986
R12342 x4.V2.n67 x4.V2.t2 20.7986
R12343 x4.V2.n68 x4.V2.t67 20.7986
R12344 x4.V2.n55 x4.V2.t49 20.7986
R12345 x4.V2.n72 x4.V2.t87 20.7986
R12346 x4.V2.n73 x4.V2.t4 20.7986
R12347 x4.V2.n74 x4.V2.t15 20.7986
R12348 x4.V2.n53 x4.V2.t80 20.7986
R12349 x4.V2.n78 x4.V2.t51 20.7986
R12350 x4.V2.n79 x4.V2.t48 20.7986
R12351 x4.V2.n80 x4.V2.t93 20.7986
R12352 x4.V2.n51 x4.V2.t78 20.7986
R12353 x4.V2.n84 x4.V2.t38 20.7986
R12354 x4.V2.n85 x4.V2.t44 20.7986
R12355 x4.V2.n86 x4.V2.t21 20.7986
R12356 x4.V2.n49 x4.V2.t50 20.7986
R12357 x4.V2.n90 x4.V2.t82 20.7986
R12358 x4.V2.n91 x4.V2.t90 20.7986
R12359 x4.V2.n92 x4.V2.t8 20.7986
R12360 x4.V2.n47 x4.V2.t46 20.7986
R12361 x4.V2.n96 x4.V2.t29 20.7986
R12362 x4.V2.n97 x4.V2.t55 20.7986
R12363 x4.V2.n98 x4.V2.t30 20.7986
R12364 x4.V2.n45 x4.V2.t91 20.7986
R12365 x4.V2.n102 x4.V2.t20 20.7986
R12366 x4.V2.n103 x4.V2.t68 20.7986
R12367 x4.V2.n104 x4.V2.t39 20.7986
R12368 x4.V2.n43 x4.V2.t66 20.7986
R12369 x4.V2.n108 x4.V2.t37 20.7986
R12370 x4.V2.n109 x4.V2.t70 20.7986
R12371 x4.V2.n110 x4.V2.t33 20.7986
R12372 x4.V2.n41 x4.V2.t65 20.7986
R12373 x4.V2.n114 x4.V2.t3 20.7986
R12374 x4.V2.n115 x4.V2.t26 20.7986
R12375 x4.V2.n116 x4.V2.t32 20.7986
R12376 x4.V2.n39 x4.V2.t1 20.7986
R12377 x4.V2.n120 x4.V2.t27 20.7986
R12378 x4.V2.n121 x4.V2.t47 20.7986
R12379 x4.V2.n122 x4.V2.t31 20.7986
R12380 x4.V2.n37 x4.V2.t69 20.7986
R12381 x4.V2.n127 x4.V2.t81 20.7986
R12382 x4.V2.n128 x4.V2.t73 20.7986
R12383 x4.V2.n35 x4.V2.t71 20.7986
R12384 x4.V2.n132 x4.V2.t72 20.7986
R12385 x4.V2.n133 x4.V2.t74 20.7986
R12386 x4.V2.n134 x4.V2.t16 20.7986
R12387 x4.V2.n33 x4.V2.t12 20.7986
R12388 x4.V2.n138 x4.V2.t57 20.7986
R12389 x4.V2.n139 x4.V2.t86 20.7986
R12390 x4.V2.n140 x4.V2.t53 20.7986
R12391 x4.V2.n31 x4.V2.t28 20.7986
R12392 x4.V2.n144 x4.V2.t58 20.7986
R12393 x4.V2.n145 x4.V2.t14 20.7986
R12394 x4.V2.n147 x4.V2.t7 20.7986
R12395 x4.V2.n146 x4.V2.t24 20.7986
R12396 x4.V2.n24 x4.V2.n23 19.9925
R12397 x4.V2.n22 x4.V2.n21 19.9925
R12398 x4.V2.n12 x4.V2.n11 19.9842
R12399 x4.V2.n10 x4.V2.n9 19.9842
R12400 x4.V2.n8 x4.V2.n7 19.9842
R12401 x4.V2.n6 x4.V2.n5 19.9842
R12402 x4.V2.n4 x4.V2.n3 19.9842
R12403 x4.V2.n2 x4.V2.n1 19.9842
R12404 x4.V2.n20 x4.V2.n19 19.9788
R12405 x4.V2.n18 x4.V2.n17 19.9788
R12406 x4.V2.n16 x4.V2.n15 19.9788
R12407 x4.V2.n14 x4.V2.n13 19.9788
R12408 x4.V2.n26 x4.V2.n25 19.0358
R12409 x4.V2.n28 x4.V2.t92 17.8929
R12410 x4.V2.n150 x4.V2.n149 15.6943
R12411 x4.V2.n151 x4.V2 12.8318
R12412 x4.V2.n59 x4.V2.t56 7.69716
R12413 x4.V2.n147 x4.V2.n146 6.93383
R12414 x4.V2.n147 x4.V2.n145 6.93383
R12415 x4.V2.n145 x4.V2.n144 6.93383
R12416 x4.V2.n144 x4.V2.n31 6.93383
R12417 x4.V2.n140 x4.V2.n31 6.93383
R12418 x4.V2.n140 x4.V2.n139 6.93383
R12419 x4.V2.n139 x4.V2.n138 6.93383
R12420 x4.V2.n138 x4.V2.n33 6.93383
R12421 x4.V2.n134 x4.V2.n33 6.93383
R12422 x4.V2.n134 x4.V2.n133 6.93383
R12423 x4.V2.n133 x4.V2.n132 6.93383
R12424 x4.V2.n132 x4.V2.n35 6.93383
R12425 x4.V2.n128 x4.V2.n35 6.93383
R12426 x4.V2.n128 x4.V2.n127 6.93383
R12427 x4.V2.n127 x4.V2.n126 6.93383
R12428 x4.V2.n126 x4.V2.n37 6.93383
R12429 x4.V2.n122 x4.V2.n37 6.93383
R12430 x4.V2.n122 x4.V2.n121 6.93383
R12431 x4.V2.n121 x4.V2.n120 6.93383
R12432 x4.V2.n120 x4.V2.n39 6.93383
R12433 x4.V2.n116 x4.V2.n39 6.93383
R12434 x4.V2.n116 x4.V2.n115 6.93383
R12435 x4.V2.n115 x4.V2.n114 6.93383
R12436 x4.V2.n114 x4.V2.n41 6.93383
R12437 x4.V2.n110 x4.V2.n41 6.93383
R12438 x4.V2.n110 x4.V2.n109 6.93383
R12439 x4.V2.n109 x4.V2.n108 6.93383
R12440 x4.V2.n108 x4.V2.n43 6.93383
R12441 x4.V2.n104 x4.V2.n43 6.93383
R12442 x4.V2.n104 x4.V2.n103 6.93383
R12443 x4.V2.n103 x4.V2.n102 6.93383
R12444 x4.V2.n102 x4.V2.n45 6.93383
R12445 x4.V2.n98 x4.V2.n45 6.93383
R12446 x4.V2.n98 x4.V2.n97 6.93383
R12447 x4.V2.n97 x4.V2.n96 6.93383
R12448 x4.V2.n96 x4.V2.n47 6.93383
R12449 x4.V2.n92 x4.V2.n47 6.93383
R12450 x4.V2.n92 x4.V2.n91 6.93383
R12451 x4.V2.n91 x4.V2.n90 6.93383
R12452 x4.V2.n90 x4.V2.n49 6.93383
R12453 x4.V2.n86 x4.V2.n49 6.93383
R12454 x4.V2.n86 x4.V2.n85 6.93383
R12455 x4.V2.n85 x4.V2.n84 6.93383
R12456 x4.V2.n84 x4.V2.n51 6.93383
R12457 x4.V2.n80 x4.V2.n51 6.93383
R12458 x4.V2.n80 x4.V2.n79 6.93383
R12459 x4.V2.n79 x4.V2.n78 6.93383
R12460 x4.V2.n78 x4.V2.n53 6.93383
R12461 x4.V2.n74 x4.V2.n53 6.93383
R12462 x4.V2.n74 x4.V2.n73 6.93383
R12463 x4.V2.n73 x4.V2.n72 6.93383
R12464 x4.V2.n72 x4.V2.n55 6.93383
R12465 x4.V2.n68 x4.V2.n55 6.93383
R12466 x4.V2.n68 x4.V2.n67 6.93383
R12467 x4.V2.n67 x4.V2.n66 6.93383
R12468 x4.V2.n66 x4.V2.n57 6.93383
R12469 x4.V2.n58 x4.V2.n57 6.93383
R12470 x4.V2.n60 x4.V2.n59 6.93383
R12471 x4.V2.n61 x4.V2.n60 6.93383
R12472 x4.V2.n62 x4.V2.n61 6.93383
R12473 x4.V2.n28 x4.V2.n27 5.42932
R12474 x4.V2.n19 x4.V2.t43 3.77447
R12475 x4.V2.n19 x4.V2.t60 3.77447
R12476 x4.V2.n17 x4.V2.t62 3.77447
R12477 x4.V2.n17 x4.V2.t42 3.77447
R12478 x4.V2.n15 x4.V2.t19 3.77447
R12479 x4.V2.n15 x4.V2.t18 3.77447
R12480 x4.V2.n13 x4.V2.t61 3.77447
R12481 x4.V2.n13 x4.V2.t17 3.77447
R12482 x4.V2.n11 x4.V2.t83 3.75732
R12483 x4.V2.n11 x4.V2.t84 3.75732
R12484 x4.V2.n9 x4.V2.t22 3.75732
R12485 x4.V2.n9 x4.V2.t23 3.75732
R12486 x4.V2.n7 x4.V2.t63 3.75732
R12487 x4.V2.n7 x4.V2.t6 3.75732
R12488 x4.V2.n5 x4.V2.t11 3.75732
R12489 x4.V2.n5 x4.V2.t10 3.75732
R12490 x4.V2.n3 x4.V2.t5 3.75732
R12491 x4.V2.n3 x4.V2.t77 3.75732
R12492 x4.V2.n1 x4.V2.t85 3.75732
R12493 x4.V2.n1 x4.V2.t9 3.75732
R12494 x4.V2.n0 x4.V2.t79 3.75732
R12495 x4.V2.n0 x4.V2.t76 3.75732
R12496 x4.V2.n23 x4.V2.t25 3.55534
R12497 x4.V2.n23 x4.V2.t35 3.55534
R12498 x4.V2.n21 x4.V2.t34 3.55534
R12499 x4.V2.n21 x4.V2.t36 3.55534
R12500 x4.V2.n25 x4.V2.t40 3.39475
R12501 x4.V2.n25 x4.V2.t41 3.39475
R12502 x4.V2.n14 x4.V2.n12 1.55606
R12503 x4.V2.n22 x4.V2.n20 1.55606
R12504 x4.V2.n26 x4.V2.n24 1.55606
R12505 x4.V2.n27 x4.V2.n26 1.55606
R12506 x4.V2.n16 x4.V2.n14 0.898069
R12507 x4.V2.n20 x4.V2.n18 0.898069
R12508 x4.V2.n4 x4.V2.n2 0.896333
R12509 x4.V2.n6 x4.V2.n4 0.896333
R12510 x4.V2.n8 x4.V2.n6 0.896333
R12511 x4.V2.n12 x4.V2.n10 0.896333
R12512 x4.V2.n24 x4.V2.n22 0.896333
R12513 x4.V2.n10 x4.V2.n8 0.894597
R12514 x4.V2.n18 x4.V2.n16 0.894597
R12515 x4.V2.n64 x4.V2.n57 0.7755
R12516 x4.V2.n66 x4.V2.n65 0.7755
R12517 x4.V2.n67 x4.V2.n56 0.7755
R12518 x4.V2.n69 x4.V2.n68 0.7755
R12519 x4.V2.n70 x4.V2.n55 0.7755
R12520 x4.V2.n72 x4.V2.n71 0.7755
R12521 x4.V2.n73 x4.V2.n54 0.7755
R12522 x4.V2.n75 x4.V2.n74 0.7755
R12523 x4.V2.n76 x4.V2.n53 0.7755
R12524 x4.V2.n78 x4.V2.n77 0.7755
R12525 x4.V2.n79 x4.V2.n52 0.7755
R12526 x4.V2.n81 x4.V2.n80 0.7755
R12527 x4.V2.n82 x4.V2.n51 0.7755
R12528 x4.V2.n84 x4.V2.n83 0.7755
R12529 x4.V2.n85 x4.V2.n50 0.7755
R12530 x4.V2.n87 x4.V2.n86 0.7755
R12531 x4.V2.n88 x4.V2.n49 0.7755
R12532 x4.V2.n90 x4.V2.n89 0.7755
R12533 x4.V2.n91 x4.V2.n48 0.7755
R12534 x4.V2.n93 x4.V2.n92 0.7755
R12535 x4.V2.n94 x4.V2.n47 0.7755
R12536 x4.V2.n96 x4.V2.n95 0.7755
R12537 x4.V2.n97 x4.V2.n46 0.7755
R12538 x4.V2.n99 x4.V2.n98 0.7755
R12539 x4.V2.n100 x4.V2.n45 0.7755
R12540 x4.V2.n102 x4.V2.n101 0.7755
R12541 x4.V2.n103 x4.V2.n44 0.7755
R12542 x4.V2.n105 x4.V2.n104 0.7755
R12543 x4.V2.n106 x4.V2.n43 0.7755
R12544 x4.V2.n108 x4.V2.n107 0.7755
R12545 x4.V2.n109 x4.V2.n42 0.7755
R12546 x4.V2.n111 x4.V2.n110 0.7755
R12547 x4.V2.n112 x4.V2.n41 0.7755
R12548 x4.V2.n114 x4.V2.n113 0.7755
R12549 x4.V2.n115 x4.V2.n40 0.7755
R12550 x4.V2.n117 x4.V2.n116 0.7755
R12551 x4.V2.n118 x4.V2.n39 0.7755
R12552 x4.V2.n120 x4.V2.n119 0.7755
R12553 x4.V2.n121 x4.V2.n38 0.7755
R12554 x4.V2.n123 x4.V2.n122 0.7755
R12555 x4.V2.n124 x4.V2.n37 0.7755
R12556 x4.V2.n127 x4.V2.n36 0.7755
R12557 x4.V2.n129 x4.V2.n128 0.7755
R12558 x4.V2.n130 x4.V2.n35 0.7755
R12559 x4.V2.n132 x4.V2.n131 0.7755
R12560 x4.V2.n133 x4.V2.n34 0.7755
R12561 x4.V2.n135 x4.V2.n134 0.7755
R12562 x4.V2.n136 x4.V2.n33 0.7755
R12563 x4.V2.n138 x4.V2.n137 0.7755
R12564 x4.V2.n139 x4.V2.n32 0.7755
R12565 x4.V2.n141 x4.V2.n140 0.7755
R12566 x4.V2.n142 x4.V2.n31 0.7755
R12567 x4.V2.n144 x4.V2.n143 0.7755
R12568 x4.V2.n145 x4.V2.n29 0.7755
R12569 x4.V2.n148 x4.V2.n147 0.7755
R12570 x4.V2.n126 x4.V2.n125 0.7755
R12571 x4.V2.n59 x4.V2.t45 0.763824
R12572 x4.V2.n60 x4.V2.t54 0.763824
R12573 x4.V2.n61 x4.V2.t88 0.763824
R12574 x4.V2.n126 x4.V2.t0 0.763824
R12575 x4.V2.n63 x4.V2.n62 0.684283
R12576 x4.V2.n63 x4.V2.n58 0.629383
R12577 x4.V2.n146 x4.V2.n30 0.629383
R12578 x4.V2 x4.V2.n28 0.558313
R12579 x4.V2.n151 x4.V2.n150 0.343208
R12580 x4.V2.n64 x4.V2.n63 0.145085
R12581 x4.V2.n148 x4.V2.n30 0.145085
R12582 x4.V2.n65 x4.V2.n64 0.0682083
R12583 x4.V2.n65 x4.V2.n56 0.0682083
R12584 x4.V2.n69 x4.V2.n56 0.0682083
R12585 x4.V2.n70 x4.V2.n69 0.0682083
R12586 x4.V2.n71 x4.V2.n70 0.0682083
R12587 x4.V2.n71 x4.V2.n54 0.0682083
R12588 x4.V2.n75 x4.V2.n54 0.0682083
R12589 x4.V2.n76 x4.V2.n75 0.0682083
R12590 x4.V2.n77 x4.V2.n76 0.0682083
R12591 x4.V2.n77 x4.V2.n52 0.0682083
R12592 x4.V2.n81 x4.V2.n52 0.0682083
R12593 x4.V2.n82 x4.V2.n81 0.0682083
R12594 x4.V2.n83 x4.V2.n82 0.0682083
R12595 x4.V2.n83 x4.V2.n50 0.0682083
R12596 x4.V2.n87 x4.V2.n50 0.0682083
R12597 x4.V2.n88 x4.V2.n87 0.0682083
R12598 x4.V2.n89 x4.V2.n88 0.0682083
R12599 x4.V2.n89 x4.V2.n48 0.0682083
R12600 x4.V2.n93 x4.V2.n48 0.0682083
R12601 x4.V2.n94 x4.V2.n93 0.0682083
R12602 x4.V2.n95 x4.V2.n94 0.0682083
R12603 x4.V2.n95 x4.V2.n46 0.0682083
R12604 x4.V2.n99 x4.V2.n46 0.0682083
R12605 x4.V2.n100 x4.V2.n99 0.0682083
R12606 x4.V2.n101 x4.V2.n100 0.0682083
R12607 x4.V2.n101 x4.V2.n44 0.0682083
R12608 x4.V2.n105 x4.V2.n44 0.0682083
R12609 x4.V2.n106 x4.V2.n105 0.0682083
R12610 x4.V2.n107 x4.V2.n106 0.0682083
R12611 x4.V2.n107 x4.V2.n42 0.0682083
R12612 x4.V2.n111 x4.V2.n42 0.0682083
R12613 x4.V2.n112 x4.V2.n111 0.0682083
R12614 x4.V2.n113 x4.V2.n112 0.0682083
R12615 x4.V2.n113 x4.V2.n40 0.0682083
R12616 x4.V2.n117 x4.V2.n40 0.0682083
R12617 x4.V2.n118 x4.V2.n117 0.0682083
R12618 x4.V2.n119 x4.V2.n118 0.0682083
R12619 x4.V2.n119 x4.V2.n38 0.0682083
R12620 x4.V2.n123 x4.V2.n38 0.0682083
R12621 x4.V2.n124 x4.V2.n123 0.0682083
R12622 x4.V2.n125 x4.V2.n124 0.0682083
R12623 x4.V2.n125 x4.V2.n36 0.0682083
R12624 x4.V2.n129 x4.V2.n36 0.0682083
R12625 x4.V2.n130 x4.V2.n129 0.0682083
R12626 x4.V2.n131 x4.V2.n130 0.0682083
R12627 x4.V2.n131 x4.V2.n34 0.0682083
R12628 x4.V2.n135 x4.V2.n34 0.0682083
R12629 x4.V2.n136 x4.V2.n135 0.0682083
R12630 x4.V2.n137 x4.V2.n136 0.0682083
R12631 x4.V2.n137 x4.V2.n32 0.0682083
R12632 x4.V2.n141 x4.V2.n32 0.0682083
R12633 x4.V2.n142 x4.V2.n141 0.0682083
R12634 x4.V2.n143 x4.V2.n142 0.0682083
R12635 x4.V2.n143 x4.V2.n29 0.0682083
R12636 x4.V2 x4.V2.n151 0.063
R12637 x4.V2.n149 x4.V2.n29 0.058081
R12638 x4.V2.n149 x4.V2.n148 0.0106273
R12639 D43v3.n7 D43v3.n6 873.303
R12640 D43v3 D43v3.n7 585
R12641 D43v3.t1 D43v3 506.99
R12642 D43v3 D43v3.t0 150.315
R12643 D43v3.n7 D43v3.t1 147.756
R12644 D43v3.n0 D43v3.t18 105.097
R12645 D43v3.n1 D43v3.t19 105.097
R12646 D43v3.n3 D43v3.t14 104.712
R12647 D43v3.n3 D43v3.t28 104.712
R12648 D43v3.n3 D43v3.t26 104.712
R12649 D43v3.n3 D43v3.t4 104.712
R12650 D43v3.n0 D43v3.t12 104.712
R12651 D43v3.n0 D43v3.t10 104.712
R12652 D43v3.n0 D43v3.t24 104.712
R12653 D43v3.n0 D43v3.t22 104.712
R12654 D43v3.n0 D43v3.t2 104.712
R12655 D43v3.n0 D43v3.t8 104.712
R12656 D43v3.n0 D43v3.t6 104.712
R12657 D43v3.n0 D43v3.t20 104.712
R12658 D43v3.n2 D43v3.t15 104.712
R12659 D43v3.n2 D43v3.t29 104.712
R12660 D43v3.n2 D43v3.t27 104.712
R12661 D43v3.n2 D43v3.t5 104.712
R12662 D43v3.n1 D43v3.t13 104.712
R12663 D43v3.n1 D43v3.t11 104.712
R12664 D43v3.n1 D43v3.t25 104.712
R12665 D43v3.n1 D43v3.t23 104.712
R12666 D43v3.n1 D43v3.t3 104.712
R12667 D43v3.n1 D43v3.t9 104.712
R12668 D43v3.n1 D43v3.t7 104.712
R12669 D43v3.n1 D43v3.t21 104.712
R12670 D43v3.n4 D43v3.t16 99.9956
R12671 D43v3.n5 D43v3.t17 99.9875
R12672 D43v3.n3 D43v3 14.5286
R12673 D43v3.n5 D43v3.n4 13.4337
R12674 D43v3 D43v3.n2 9.62237
R12675 D43v3.n6 D43v3 4.99562
R12676 D43v3.n2 D43v3.n1 4.838
R12677 D43v3.n3 D43v3.n0 4.838
R12678 D43v3.n2 D43v3.n5 4.72499
R12679 D43v3.n4 D43v3.n3 4.71691
R12680 D43v3 D43v3.n6 2.70619
R12681 a_6164_n9984.n1 a_6164_n9984.t10 24.2469
R12682 a_6164_n9984.n26 a_6164_n9984.t23 21.6428
R12683 a_6164_n9984.n26 a_6164_n9984.t26 21.5736
R12684 a_6164_n9984.n25 a_6164_n9984.t21 21.5736
R12685 a_6164_n9984.n24 a_6164_n9984.t28 21.5736
R12686 a_6164_n9984.n23 a_6164_n9984.t29 21.5736
R12687 a_6164_n9984.n22 a_6164_n9984.t24 21.5736
R12688 a_6164_n9984.n21 a_6164_n9984.t19 21.5736
R12689 a_6164_n9984.n20 a_6164_n9984.t22 21.5736
R12690 a_6164_n9984.n19 a_6164_n9984.t18 21.5736
R12691 a_6164_n9984.n18 a_6164_n9984.t2 21.5736
R12692 a_6164_n9984.n17 a_6164_n9984.t3 21.5736
R12693 a_6164_n9984.n16 a_6164_n9984.t1 21.5736
R12694 a_6164_n9984.n15 a_6164_n9984.t25 21.5736
R12695 a_6164_n9984.n14 a_6164_n9984.t20 21.5736
R12696 a_6164_n9984.n13 a_6164_n9984.t27 21.5736
R12697 a_6164_n9984.n1 a_6164_n9984.n0 19.6822
R12698 a_6164_n9984.n3 a_6164_n9984.n2 19.6822
R12699 a_6164_n9984.n5 a_6164_n9984.n4 19.6822
R12700 a_6164_n9984.n7 a_6164_n9984.n6 19.6822
R12701 a_6164_n9984.n9 a_6164_n9984.n8 19.6822
R12702 a_6164_n9984.n11 a_6164_n9984.n10 19.6822
R12703 a_6164_n9984.n12 a_6164_n9984.t9 18.7631
R12704 a_6164_n9984.n0 a_6164_n9984.t4 3.75732
R12705 a_6164_n9984.n0 a_6164_n9984.t11 3.75732
R12706 a_6164_n9984.n2 a_6164_n9984.t16 3.75732
R12707 a_6164_n9984.n2 a_6164_n9984.t5 3.75732
R12708 a_6164_n9984.n4 a_6164_n9984.t13 3.75732
R12709 a_6164_n9984.n4 a_6164_n9984.t12 3.75732
R12710 a_6164_n9984.n6 a_6164_n9984.t7 3.75732
R12711 a_6164_n9984.n6 a_6164_n9984.t6 3.75732
R12712 a_6164_n9984.n8 a_6164_n9984.t14 3.75732
R12713 a_6164_n9984.n8 a_6164_n9984.t17 3.75732
R12714 a_6164_n9984.n10 a_6164_n9984.t8 3.75732
R12715 a_6164_n9984.n10 a_6164_n9984.t15 3.75732
R12716 a_6164_n9984.n12 a_6164_n9984.n11 3.21198
R12717 a_6164_n9984.t0 a_6164_n9984.n27 1.53882
R12718 a_6164_n9984.n13 a_6164_n9984.n12 0.943131
R12719 a_6164_n9984.n11 a_6164_n9984.n9 0.808313
R12720 a_6164_n9984.n9 a_6164_n9984.n7 0.80675
R12721 a_6164_n9984.n7 a_6164_n9984.n5 0.80675
R12722 a_6164_n9984.n5 a_6164_n9984.n3 0.80675
R12723 a_6164_n9984.n3 a_6164_n9984.n1 0.80675
R12724 a_6164_n9984.n14 a_6164_n9984.n13 0.0696489
R12725 a_6164_n9984.n15 a_6164_n9984.n14 0.0696489
R12726 a_6164_n9984.n16 a_6164_n9984.n15 0.0696489
R12727 a_6164_n9984.n17 a_6164_n9984.n16 0.0696489
R12728 a_6164_n9984.n18 a_6164_n9984.n17 0.0696489
R12729 a_6164_n9984.n19 a_6164_n9984.n18 0.0696489
R12730 a_6164_n9984.n20 a_6164_n9984.n19 0.0696489
R12731 a_6164_n9984.n21 a_6164_n9984.n20 0.0696489
R12732 a_6164_n9984.n22 a_6164_n9984.n21 0.0696489
R12733 a_6164_n9984.n23 a_6164_n9984.n22 0.0696489
R12734 a_6164_n9984.n24 a_6164_n9984.n23 0.0696489
R12735 a_6164_n9984.n25 a_6164_n9984.n24 0.0696489
R12736 a_6164_n9984.n27 a_6164_n9984.n25 0.0696489
R12737 a_6164_n9984.n27 a_6164_n9984.n26 0.0696489
R12738 AVOUT2.n0 AVOUT2.t38 491.555
R12739 AVOUT2.n6 AVOUT2.t27 25.5864
R12740 AVOUT2.n8 AVOUT2.t32 21.5504
R12741 AVOUT2.n8 AVOUT2.t17 21.4809
R12742 AVOUT2.n9 AVOUT2.t29 21.4809
R12743 AVOUT2.n10 AVOUT2.t3 21.4809
R12744 AVOUT2.n11 AVOUT2.t10 21.4809
R12745 AVOUT2.n12 AVOUT2.t9 21.4809
R12746 AVOUT2.n13 AVOUT2.t12 21.4809
R12747 AVOUT2.n14 AVOUT2.t20 21.4809
R12748 AVOUT2.n15 AVOUT2.t13 21.4809
R12749 AVOUT2.n16 AVOUT2.t26 21.4809
R12750 AVOUT2.n17 AVOUT2.t35 21.4809
R12751 AVOUT2.n18 AVOUT2.t33 21.4809
R12752 AVOUT2.n19 AVOUT2.t18 21.4809
R12753 AVOUT2.n20 AVOUT2.t0 21.4809
R12754 AVOUT2.n21 AVOUT2.t31 21.4809
R12755 AVOUT2.n22 AVOUT2.t25 21.4809
R12756 AVOUT2.n24 AVOUT2.t16 21.4809
R12757 AVOUT2.n25 AVOUT2.t21 21.4809
R12758 AVOUT2.n26 AVOUT2.t36 21.4809
R12759 AVOUT2.n27 AVOUT2.t22 21.4809
R12760 AVOUT2.n28 AVOUT2.t8 21.4809
R12761 AVOUT2.n29 AVOUT2.t2 21.4809
R12762 AVOUT2.n30 AVOUT2.t1 21.4809
R12763 AVOUT2.n31 AVOUT2.t34 21.4809
R12764 AVOUT2.n32 AVOUT2.t7 21.4809
R12765 AVOUT2.n33 AVOUT2.t14 21.4809
R12766 AVOUT2.n34 AVOUT2.t37 21.4809
R12767 AVOUT2.n35 AVOUT2.t28 21.4809
R12768 AVOUT2.n36 AVOUT2.t30 21.4809
R12769 AVOUT2.n37 AVOUT2.t11 21.4809
R12770 AVOUT2.n38 AVOUT2.t19 21.4809
R12771 AVOUT2.n39 AVOUT2.t15 21.4809
R12772 AVOUT2.n3 AVOUT2.n1 13.4669
R12773 AVOUT2.n3 AVOUT2.n2 13.3799
R12774 AVOUT2.n7 AVOUT2.n0 9.895
R12775 AVOUT2.n23 AVOUT2.n7 8.01275
R12776 AVOUT2.n40 AVOUT2 5.14269
R12777 AVOUT2.n5 AVOUT2.t6 4.35292
R12778 AVOUT2.n6 AVOUT2.n5 3.83074
R12779 AVOUT2.n5 AVOUT2.n4 3.24934
R12780 AVOUT2.n4 AVOUT2 2.58592
R12781 AVOUT2.n4 AVOUT2.n3 2.00817
R12782 AVOUT2.n1 AVOUT2.t5 1.45813
R12783 AVOUT2.n1 AVOUT2.t24 1.45813
R12784 AVOUT2.n2 AVOUT2.t23 1.45813
R12785 AVOUT2.n2 AVOUT2.t4 1.45813
R12786 AVOUT2.n0 AVOUT2 1.34958
R12787 AVOUT2.n40 AVOUT2.n39 0.633643
R12788 AVOUT2.n32 AVOUT2.n31 0.223778
R12789 AVOUT2.n36 AVOUT2.n35 0.205963
R12790 AVOUT2.n38 AVOUT2.n37 0.188148
R12791 AVOUT2.n39 AVOUT2.n38 0.15727
R12792 AVOUT2.n7 AVOUT2.n6 0.14011
R12793 AVOUT2.n24 AVOUT2.n23 0.138564
R12794 AVOUT2.n9 AVOUT2.n8 0.0699774
R12795 AVOUT2.n10 AVOUT2.n9 0.0699774
R12796 AVOUT2.n11 AVOUT2.n10 0.0699774
R12797 AVOUT2.n12 AVOUT2.n11 0.0699774
R12798 AVOUT2.n13 AVOUT2.n12 0.0699774
R12799 AVOUT2.n14 AVOUT2.n13 0.0699774
R12800 AVOUT2.n15 AVOUT2.n14 0.0699774
R12801 AVOUT2.n16 AVOUT2.n15 0.0699774
R12802 AVOUT2.n17 AVOUT2.n16 0.0699774
R12803 AVOUT2.n18 AVOUT2.n17 0.0699774
R12804 AVOUT2.n19 AVOUT2.n18 0.0699774
R12805 AVOUT2.n20 AVOUT2.n19 0.0699774
R12806 AVOUT2.n21 AVOUT2.n20 0.0699774
R12807 AVOUT2.n22 AVOUT2.n21 0.0699774
R12808 AVOUT2.n25 AVOUT2.n24 0.0699774
R12809 AVOUT2.n26 AVOUT2.n25 0.0699774
R12810 AVOUT2.n27 AVOUT2.n26 0.0699774
R12811 AVOUT2.n28 AVOUT2.n27 0.0699774
R12812 AVOUT2.n29 AVOUT2.n28 0.0699774
R12813 AVOUT2.n30 AVOUT2.n29 0.0699774
R12814 AVOUT2.n31 AVOUT2.n30 0.0699774
R12815 AVOUT2.n33 AVOUT2.n32 0.0699774
R12816 AVOUT2.n34 AVOUT2.n33 0.0699774
R12817 AVOUT2.n35 AVOUT2.n34 0.0699774
R12818 AVOUT2.n37 AVOUT2.n36 0.0699774
R12819 AVOUT2 AVOUT2.n40 0.063
R12820 AVOUT2.n23 AVOUT2.n22 0.0583979
R12821 D33v3.n5 D33v3.n4 873.303
R12822 D33v3 D33v3.n5 585
R12823 D33v3.t1 D33v3 506.99
R12824 D33v3 D33v3.t0 150.315
R12825 D33v3.n5 D33v3.t1 147.756
R12826 D33v3.n0 D33v3.t4 104.861
R12827 D33v3.n1 D33v3.t5 104.861
R12828 D33v3.n0 D33v3.t10 104.469
R12829 D33v3.n0 D33v3.t8 104.469
R12830 D33v3.n0 D33v3.t12 104.469
R12831 D33v3.n0 D33v3.t14 104.469
R12832 D33v3.n0 D33v3.t16 104.469
R12833 D33v3.n0 D33v3.t6 104.469
R12834 D33v3.n1 D33v3.t11 104.469
R12835 D33v3.n1 D33v3.t9 104.469
R12836 D33v3.n1 D33v3.t13 104.469
R12837 D33v3.n1 D33v3.t15 104.469
R12838 D33v3.n1 D33v3.t17 104.469
R12839 D33v3.n1 D33v3.t7 104.469
R12840 D33v3.n2 D33v3.t2 99.8073
R12841 D33v3.n3 D33v3.t3 99.6942
R12842 D33v3.n3 D33v3.n2 13.4361
R12843 D33v3.n0 D33v3 10.7114
R12844 D33v3.n1 D33v3.n3 7.19034
R12845 D33v3.n2 D33v3.n0 7.0772
R12846 D33v3 D33v3.n1 5.80519
R12847 D33v3.n4 D33v3 4.99562
R12848 D33v3 D33v3.n4 2.70619
R12849 a_3720_n9984.n1 a_3720_n9984.t10 24.2695
R12850 a_3720_n9984.n13 a_3720_n9984.t14 21.6429
R12851 a_3720_n9984.n12 a_3720_n9984.t1 21.5736
R12852 a_3720_n9984.n11 a_3720_n9984.t2 21.5736
R12853 a_3720_n9984.n10 a_3720_n9984.t13 21.5736
R12854 a_3720_n9984.n9 a_3720_n9984.t15 21.5736
R12855 a_3720_n9984.n8 a_3720_n9984.t12 21.5736
R12856 a_3720_n9984.n7 a_3720_n9984.t11 21.5736
R12857 a_3720_n9984.n1 a_3720_n9984.n0 19.6768
R12858 a_3720_n9984.n3 a_3720_n9984.n2 19.6768
R12859 a_3720_n9984.n5 a_3720_n9984.n4 19.6768
R12860 a_3720_n9984.n6 a_3720_n9984.t9 18.7802
R12861 a_3720_n9984.n6 a_3720_n9984.n5 5.44609
R12862 a_3720_n9984.n0 a_3720_n9984.t7 3.77447
R12863 a_3720_n9984.n0 a_3720_n9984.t6 3.77447
R12864 a_3720_n9984.n2 a_3720_n9984.t4 3.77447
R12865 a_3720_n9984.n2 a_3720_n9984.t5 3.77447
R12866 a_3720_n9984.n4 a_3720_n9984.t8 3.77447
R12867 a_3720_n9984.n4 a_3720_n9984.t3 3.77447
R12868 a_3720_n9984.t0 a_3720_n9984.n13 1.53882
R12869 a_3720_n9984.n7 a_3720_n9984.n6 1.07925
R12870 a_3720_n9984.n5 a_3720_n9984.n3 0.808313
R12871 a_3720_n9984.n3 a_3720_n9984.n1 0.808313
R12872 a_3720_n9984.n8 a_3720_n9984.n7 0.0698128
R12873 a_3720_n9984.n9 a_3720_n9984.n8 0.0698128
R12874 a_3720_n9984.n10 a_3720_n9984.n9 0.0698128
R12875 a_3720_n9984.n11 a_3720_n9984.n10 0.0698128
R12876 a_3720_n9984.n12 a_3720_n9984.n11 0.0698128
R12877 a_3720_n9984.n13 a_3720_n9984.n12 0.0698128
R12878 a_6164_n4916.n1 a_6164_n4916.t11 24.2469
R12879 a_6164_n4916.n14 a_6164_n4916.t29 21.6428
R12880 a_6164_n4916.n14 a_6164_n4916.t28 21.5736
R12881 a_6164_n4916.n15 a_6164_n4916.t19 21.5736
R12882 a_6164_n4916.n16 a_6164_n4916.t2 21.5736
R12883 a_6164_n4916.n17 a_6164_n4916.t3 21.5736
R12884 a_6164_n4916.n18 a_6164_n4916.t26 21.5736
R12885 a_6164_n4916.n19 a_6164_n4916.t1 21.5736
R12886 a_6164_n4916.n20 a_6164_n4916.t4 21.5736
R12887 a_6164_n4916.n21 a_6164_n4916.t24 21.5736
R12888 a_6164_n4916.n22 a_6164_n4916.t20 21.5736
R12889 a_6164_n4916.n23 a_6164_n4916.t21 21.5736
R12890 a_6164_n4916.n24 a_6164_n4916.t25 21.5736
R12891 a_6164_n4916.n25 a_6164_n4916.t23 21.5736
R12892 a_6164_n4916.n26 a_6164_n4916.t27 21.5736
R12893 a_6164_n4916.n13 a_6164_n4916.t22 21.5736
R12894 a_6164_n4916.n1 a_6164_n4916.n0 19.6822
R12895 a_6164_n4916.n3 a_6164_n4916.n2 19.6822
R12896 a_6164_n4916.n5 a_6164_n4916.n4 19.6822
R12897 a_6164_n4916.n7 a_6164_n4916.n6 19.6822
R12898 a_6164_n4916.n9 a_6164_n4916.n8 19.6822
R12899 a_6164_n4916.n11 a_6164_n4916.n10 19.6822
R12900 a_6164_n4916.n12 a_6164_n4916.t10 18.7631
R12901 a_6164_n4916.n0 a_6164_n4916.t5 3.75732
R12902 a_6164_n4916.n0 a_6164_n4916.t12 3.75732
R12903 a_6164_n4916.n2 a_6164_n4916.t17 3.75732
R12904 a_6164_n4916.n2 a_6164_n4916.t6 3.75732
R12905 a_6164_n4916.n4 a_6164_n4916.t14 3.75732
R12906 a_6164_n4916.n4 a_6164_n4916.t13 3.75732
R12907 a_6164_n4916.n6 a_6164_n4916.t8 3.75732
R12908 a_6164_n4916.n6 a_6164_n4916.t7 3.75732
R12909 a_6164_n4916.n8 a_6164_n4916.t15 3.75732
R12910 a_6164_n4916.n8 a_6164_n4916.t18 3.75732
R12911 a_6164_n4916.n10 a_6164_n4916.t9 3.75732
R12912 a_6164_n4916.n10 a_6164_n4916.t16 3.75732
R12913 a_6164_n4916.n12 a_6164_n4916.n11 3.21198
R12914 a_6164_n4916.t0 a_6164_n4916.n27 1.53882
R12915 a_6164_n4916.n13 a_6164_n4916.n12 0.943131
R12916 a_6164_n4916.n11 a_6164_n4916.n9 0.808313
R12917 a_6164_n4916.n9 a_6164_n4916.n7 0.80675
R12918 a_6164_n4916.n7 a_6164_n4916.n5 0.80675
R12919 a_6164_n4916.n5 a_6164_n4916.n3 0.80675
R12920 a_6164_n4916.n3 a_6164_n4916.n1 0.80675
R12921 a_6164_n4916.n27 a_6164_n4916.n13 0.0696489
R12922 a_6164_n4916.n27 a_6164_n4916.n26 0.0696489
R12923 a_6164_n4916.n26 a_6164_n4916.n25 0.0696489
R12924 a_6164_n4916.n25 a_6164_n4916.n24 0.0696489
R12925 a_6164_n4916.n24 a_6164_n4916.n23 0.0696489
R12926 a_6164_n4916.n23 a_6164_n4916.n22 0.0696489
R12927 a_6164_n4916.n22 a_6164_n4916.n21 0.0696489
R12928 a_6164_n4916.n21 a_6164_n4916.n20 0.0696489
R12929 a_6164_n4916.n20 a_6164_n4916.n19 0.0696489
R12930 a_6164_n4916.n19 a_6164_n4916.n18 0.0696489
R12931 a_6164_n4916.n18 a_6164_n4916.n17 0.0696489
R12932 a_6164_n4916.n17 a_6164_n4916.n16 0.0696489
R12933 a_6164_n4916.n16 a_6164_n4916.n15 0.0696489
R12934 a_6164_n4916.n15 a_6164_n4916.n14 0.0696489
R12935 AVOUT1.n3 AVOUT1.t38 491.555
R12936 AVOUT1.n20 AVOUT1.t11 21.4969
R12937 AVOUT1.n4 AVOUT1.t22 21.4809
R12938 AVOUT1.n5 AVOUT1.t0 21.4809
R12939 AVOUT1.n6 AVOUT1.t32 21.4809
R12940 AVOUT1.n7 AVOUT1.t25 21.4809
R12941 AVOUT1.n8 AVOUT1.t28 21.4809
R12942 AVOUT1.n9 AVOUT1.t21 21.4809
R12943 AVOUT1.n10 AVOUT1.t18 21.4809
R12944 AVOUT1.n11 AVOUT1.t26 21.4809
R12945 AVOUT1.n12 AVOUT1.t8 21.4809
R12946 AVOUT1.n13 AVOUT1.t1 21.4809
R12947 AVOUT1.n14 AVOUT1.t29 21.4809
R12948 AVOUT1.n15 AVOUT1.t4 21.4809
R12949 AVOUT1.n16 AVOUT1.t2 21.4809
R12950 AVOUT1.n17 AVOUT1.t17 21.4809
R12951 AVOUT1.n18 AVOUT1.t33 21.4809
R12952 AVOUT1.n21 AVOUT1.t35 21.4809
R12953 AVOUT1.n22 AVOUT1.t15 21.4809
R12954 AVOUT1.n23 AVOUT1.t34 21.4809
R12955 AVOUT1.n24 AVOUT1.t20 21.4809
R12956 AVOUT1.n25 AVOUT1.t19 21.4809
R12957 AVOUT1.n27 AVOUT1.t16 21.4809
R12958 AVOUT1.n28 AVOUT1.t9 21.4809
R12959 AVOUT1.n29 AVOUT1.t24 21.4809
R12960 AVOUT1.n30 AVOUT1.t3 21.4809
R12961 AVOUT1.n31 AVOUT1.t10 21.4809
R12962 AVOUT1.n32 AVOUT1.t36 21.4809
R12963 AVOUT1.n33 AVOUT1.t14 21.4809
R12964 AVOUT1.n34 AVOUT1.t31 21.4809
R12965 AVOUT1.n35 AVOUT1.t37 21.4809
R12966 AVOUT1.n36 AVOUT1.t5 21.4809
R12967 AVOUT1.n37 AVOUT1.t30 21.4809
R12968 AVOUT1.n38 AVOUT1.t23 21.4809
R12969 AVOUT1.n2 AVOUT1.n0 13.4669
R12970 AVOUT1.n2 AVOUT1.n1 13.3799
R12971 AVOUT1.n41 AVOUT1.n40 8.69177
R12972 AVOUT1.n4 AVOUT1.n3 5.19222
R12973 AVOUT1.n40 AVOUT1.n39 4.5005
R12974 AVOUT1.n43 AVOUT1.t27 4.35292
R12975 AVOUT1.n44 AVOUT1.n43 3.22372
R12976 AVOUT1.n42 AVOUT1.n41 2.91854
R12977 AVOUT1 AVOUT1.n44 2.58592
R12978 AVOUT1.n44 AVOUT1.n2 2.00817
R12979 AVOUT1.n0 AVOUT1.t6 1.45813
R12980 AVOUT1.n0 AVOUT1.t7 1.45813
R12981 AVOUT1.n1 AVOUT1.t12 1.45813
R12982 AVOUT1.n1 AVOUT1.t13 1.45813
R12983 AVOUT1.n43 AVOUT1.n42 1.45117
R12984 AVOUT1.n3 AVOUT1 1.35154
R12985 AVOUT1.n41 AVOUT1.n20 1.05966
R12986 AVOUT1.n42 AVOUT1.n19 0.642263
R12987 AVOUT1.n39 AVOUT1.n38 0.633643
R12988 AVOUT1.n40 AVOUT1 0.627062
R12989 AVOUT1.n26 AVOUT1.n20 0.562735
R12990 AVOUT1.n31 AVOUT1.n30 0.223778
R12991 AVOUT1.n35 AVOUT1.n34 0.205963
R12992 AVOUT1.n22 AVOUT1.n21 0.196462
R12993 AVOUT1.n37 AVOUT1.n36 0.188148
R12994 AVOUT1.n38 AVOUT1.n37 0.15727
R12995 AVOUT1.n5 AVOUT1.n4 0.0699774
R12996 AVOUT1.n6 AVOUT1.n5 0.0699774
R12997 AVOUT1.n7 AVOUT1.n6 0.0699774
R12998 AVOUT1.n8 AVOUT1.n7 0.0699774
R12999 AVOUT1.n9 AVOUT1.n8 0.0699774
R13000 AVOUT1.n10 AVOUT1.n9 0.0699774
R13001 AVOUT1.n11 AVOUT1.n10 0.0699774
R13002 AVOUT1.n12 AVOUT1.n11 0.0699774
R13003 AVOUT1.n13 AVOUT1.n12 0.0699774
R13004 AVOUT1.n14 AVOUT1.n13 0.0699774
R13005 AVOUT1.n15 AVOUT1.n14 0.0699774
R13006 AVOUT1.n16 AVOUT1.n15 0.0699774
R13007 AVOUT1.n17 AVOUT1.n16 0.0699774
R13008 AVOUT1.n18 AVOUT1.n17 0.0699774
R13009 AVOUT1.n23 AVOUT1.n22 0.0699774
R13010 AVOUT1.n24 AVOUT1.n23 0.0699774
R13011 AVOUT1.n25 AVOUT1.n24 0.0699774
R13012 AVOUT1.n28 AVOUT1.n27 0.0699774
R13013 AVOUT1.n29 AVOUT1.n28 0.0699774
R13014 AVOUT1.n30 AVOUT1.n29 0.0699774
R13015 AVOUT1.n32 AVOUT1.n31 0.0699774
R13016 AVOUT1.n33 AVOUT1.n32 0.0699774
R13017 AVOUT1.n34 AVOUT1.n33 0.0699774
R13018 AVOUT1.n36 AVOUT1.n35 0.0699774
R13019 AVOUT1.n39 AVOUT1 0.063
R13020 AVOUT1.n19 AVOUT1.n18 0.0610701
R13021 AVOUT1.n27 AVOUT1.n26 0.0480059
R13022 AVOUT1.n26 AVOUT1.n25 0.0224715
R13023 AVOUT1.n21 AVOUT1.n19 0.00940736
R13024 D73v3.n5 D73v3.n4 873.303
R13025 D73v3 D73v3.n5 585
R13026 D73v3.t1 D73v3 506.99
R13027 D73v3 D73v3.t0 150.315
R13028 D73v3.n5 D73v3.t1 147.756
R13029 D73v3.n0 D73v3.t9 108.13
R13030 D73v3.n1 D73v3.t8 108.13
R13031 D73v3.n0 D73v3.t5 107.737
R13032 D73v3.n0 D73v3.t7 107.737
R13033 D73v3.n1 D73v3.t2 107.737
R13034 D73v3.n1 D73v3.t4 107.737
R13035 D73v3.n1 D73v3.t6 107.737
R13036 D73v3.n2 D73v3.t3 102.909
R13037 D73v3 D73v3.n3 24.2833
R13038 D73v3.n0 D73v3 8.5005
R13039 D73v3.n1 D73v3 8.39112
R13040 D73v3.n3 D73v3.n2 6.67917
R13041 D73v3.n2 D73v3.n0 5.63477
R13042 D73v3.n4 D73v3 4.99562
R13043 D73v3.n3 D73v3.n1 3.07935
R13044 D73v3 D73v3.n4 2.70619
R13045 a_12405_n9984.n1 a_12405_n9984.t5 24.0657
R13046 a_12405_n9984.n4 a_12405_n9984.t6 21.6429
R13047 a_12405_n9984.n4 a_12405_n9984.t7 21.5736
R13048 a_12405_n9984.n3 a_12405_n9984.t1 21.5736
R13049 a_12405_n9984.n1 a_12405_n9984.n0 19.6936
R13050 a_12405_n9984.n2 a_12405_n9984.t2 18.5015
R13051 a_12405_n9984.n2 a_12405_n9984.n1 5.46945
R13052 a_12405_n9984.n0 a_12405_n9984.t3 3.55534
R13053 a_12405_n9984.n0 a_12405_n9984.t4 3.55534
R13054 a_12405_n9984.t0 a_12405_n9984.n5 1.53882
R13055 a_12405_n9984.n3 a_12405_n9984.n2 1.04507
R13056 a_12405_n9984.n5 a_12405_n9984.n3 0.0698128
R13057 a_12405_n9984.n5 a_12405_n9984.n4 0.0698128
R13058 a_3720_n4916.n1 a_3720_n4916.t9 24.2695
R13059 a_3720_n4916.n13 a_3720_n4916.t14 21.5736
R13060 a_3720_n4916.n12 a_3720_n4916.t1 21.5736
R13061 a_3720_n4916.n11 a_3720_n4916.t11 21.5736
R13062 a_3720_n4916.n10 a_3720_n4916.t12 21.5736
R13063 a_3720_n4916.n9 a_3720_n4916.t13 21.5736
R13064 a_3720_n4916.n8 a_3720_n4916.t15 21.5736
R13065 a_3720_n4916.n7 a_3720_n4916.t10 21.5736
R13066 a_3720_n4916.n1 a_3720_n4916.n0 19.6768
R13067 a_3720_n4916.n3 a_3720_n4916.n2 19.6768
R13068 a_3720_n4916.n5 a_3720_n4916.n4 19.6768
R13069 a_3720_n4916.n6 a_3720_n4916.t8 18.7802
R13070 a_3720_n4916.n6 a_3720_n4916.n5 5.44609
R13071 a_3720_n4916.n0 a_3720_n4916.t6 3.77447
R13072 a_3720_n4916.n0 a_3720_n4916.t5 3.77447
R13073 a_3720_n4916.n2 a_3720_n4916.t3 3.77447
R13074 a_3720_n4916.n2 a_3720_n4916.t4 3.77447
R13075 a_3720_n4916.n4 a_3720_n4916.t7 3.77447
R13076 a_3720_n4916.n4 a_3720_n4916.t2 3.77447
R13077 a_3720_n4916.t0 a_3720_n4916.n13 1.60814
R13078 a_3720_n4916.n7 a_3720_n4916.n6 1.07925
R13079 a_3720_n4916.n5 a_3720_n4916.n3 0.808313
R13080 a_3720_n4916.n3 a_3720_n4916.n1 0.808313
R13081 a_3720_n4916.n8 a_3720_n4916.n7 0.0698128
R13082 a_3720_n4916.n9 a_3720_n4916.n8 0.0698128
R13083 a_3720_n4916.n10 a_3720_n4916.n9 0.0698128
R13084 a_3720_n4916.n11 a_3720_n4916.n10 0.0698128
R13085 a_3720_n4916.n12 a_3720_n4916.n11 0.0698128
R13086 a_3720_n4916.n13 a_3720_n4916.n12 0.0698128
R13087 x8.V2.n130 x8.V2.t70 491.705
R13088 x8.V2.n128 x8.V2.t32 39.1599
R13089 x8.V2.n69 x8.V2.t53 21.4824
R13090 x8.V2.n18 x8.V2.t26 20.7986
R13091 x8.V2.n14 x8.V2.t24 20.7986
R13092 x8.V2.n21 x8.V2.t13 20.7986
R13093 x8.V2.n22 x8.V2.t36 20.7986
R13094 x8.V2.n12 x8.V2.t44 20.7986
R13095 x8.V2.n27 x8.V2.t55 20.7986
R13096 x8.V2.n28 x8.V2.t67 20.7986
R13097 x8.V2.n29 x8.V2.t60 20.7986
R13098 x8.V2.n10 x8.V2.t10 20.7986
R13099 x8.V2.n33 x8.V2.t12 20.7986
R13100 x8.V2.n34 x8.V2.t49 20.7986
R13101 x8.V2.n35 x8.V2.t25 20.7986
R13102 x8.V2.n8 x8.V2.t2 20.7986
R13103 x8.V2.n39 x8.V2.t9 20.7986
R13104 x8.V2.n40 x8.V2.t56 20.7986
R13105 x8.V2.n41 x8.V2.t29 20.7986
R13106 x8.V2.n6 x8.V2.t23 20.7986
R13107 x8.V2.n45 x8.V2.t50 20.7986
R13108 x8.V2.n46 x8.V2.t3 20.7986
R13109 x8.V2.n47 x8.V2.t52 20.7986
R13110 x8.V2.n4 x8.V2.t62 20.7986
R13111 x8.V2.n51 x8.V2.t17 20.7986
R13112 x8.V2.n52 x8.V2.t41 20.7986
R13113 x8.V2.n120 x8.V2.t63 20.7986
R13114 x8.V2.n119 x8.V2.t40 20.7986
R13115 x8.V2.n118 x8.V2.t11 20.7986
R13116 x8.V2.n53 x8.V2.t21 20.7986
R13117 x8.V2.n114 x8.V2.t43 20.7986
R13118 x8.V2.n113 x8.V2.t5 20.7986
R13119 x8.V2.n112 x8.V2.t65 20.7986
R13120 x8.V2.n55 x8.V2.t38 20.7986
R13121 x8.V2.n108 x8.V2.t7 20.7986
R13122 x8.V2.n107 x8.V2.t58 20.7986
R13123 x8.V2.n106 x8.V2.t6 20.7986
R13124 x8.V2.n57 x8.V2.t57 20.7986
R13125 x8.V2.n102 x8.V2.t47 20.7986
R13126 x8.V2.n101 x8.V2.t66 20.7986
R13127 x8.V2.n100 x8.V2.t39 20.7986
R13128 x8.V2.n59 x8.V2.t68 20.7986
R13129 x8.V2.n96 x8.V2.t1 20.7986
R13130 x8.V2.n95 x8.V2.t19 20.7986
R13131 x8.V2.n94 x8.V2.t54 20.7986
R13132 x8.V2.n61 x8.V2.t28 20.7986
R13133 x8.V2.n90 x8.V2.t15 20.7986
R13134 x8.V2.n89 x8.V2.t64 20.7986
R13135 x8.V2.n88 x8.V2.t61 20.7986
R13136 x8.V2.n63 x8.V2.t14 20.7986
R13137 x8.V2.n84 x8.V2.t4 20.7986
R13138 x8.V2.n83 x8.V2.t27 20.7986
R13139 x8.V2.n82 x8.V2.t22 20.7986
R13140 x8.V2.n65 x8.V2.t18 20.7986
R13141 x8.V2.n78 x8.V2.t37 20.7986
R13142 x8.V2.n77 x8.V2.t51 20.7986
R13143 x8.V2.n76 x8.V2.t16 20.7986
R13144 x8.V2.n67 x8.V2.t8 20.7986
R13145 x8.V2.n72 x8.V2.t69 20.7986
R13146 x8.V2.n71 x8.V2.t42 20.7986
R13147 x8.V2.n70 x8.V2.t48 20.7986
R13148 x8.V2.n125 x8.V2.n124 10.6258
R13149 x8.V2.n1 x8.V2.n0 10.6258
R13150 x8.V2.n15 x8.V2.t20 7.69716
R13151 x8.V2.n71 x8.V2.n70 6.93383
R13152 x8.V2.n72 x8.V2.n71 6.93383
R13153 x8.V2.n72 x8.V2.n67 6.93383
R13154 x8.V2.n76 x8.V2.n67 6.93383
R13155 x8.V2.n77 x8.V2.n76 6.93383
R13156 x8.V2.n78 x8.V2.n77 6.93383
R13157 x8.V2.n78 x8.V2.n65 6.93383
R13158 x8.V2.n82 x8.V2.n65 6.93383
R13159 x8.V2.n83 x8.V2.n82 6.93383
R13160 x8.V2.n84 x8.V2.n83 6.93383
R13161 x8.V2.n84 x8.V2.n63 6.93383
R13162 x8.V2.n88 x8.V2.n63 6.93383
R13163 x8.V2.n89 x8.V2.n88 6.93383
R13164 x8.V2.n90 x8.V2.n89 6.93383
R13165 x8.V2.n90 x8.V2.n61 6.93383
R13166 x8.V2.n94 x8.V2.n61 6.93383
R13167 x8.V2.n95 x8.V2.n94 6.93383
R13168 x8.V2.n96 x8.V2.n95 6.93383
R13169 x8.V2.n96 x8.V2.n59 6.93383
R13170 x8.V2.n100 x8.V2.n59 6.93383
R13171 x8.V2.n101 x8.V2.n100 6.93383
R13172 x8.V2.n102 x8.V2.n101 6.93383
R13173 x8.V2.n102 x8.V2.n57 6.93383
R13174 x8.V2.n106 x8.V2.n57 6.93383
R13175 x8.V2.n107 x8.V2.n106 6.93383
R13176 x8.V2.n108 x8.V2.n107 6.93383
R13177 x8.V2.n108 x8.V2.n55 6.93383
R13178 x8.V2.n112 x8.V2.n55 6.93383
R13179 x8.V2.n113 x8.V2.n112 6.93383
R13180 x8.V2.n114 x8.V2.n113 6.93383
R13181 x8.V2.n114 x8.V2.n53 6.93383
R13182 x8.V2.n118 x8.V2.n53 6.93383
R13183 x8.V2.n119 x8.V2.n118 6.93383
R13184 x8.V2.n120 x8.V2.n119 6.93383
R13185 x8.V2.n120 x8.V2.n52 6.93383
R13186 x8.V2.n52 x8.V2.n51 6.93383
R13187 x8.V2.n51 x8.V2.n4 6.93383
R13188 x8.V2.n47 x8.V2.n4 6.93383
R13189 x8.V2.n47 x8.V2.n46 6.93383
R13190 x8.V2.n46 x8.V2.n45 6.93383
R13191 x8.V2.n45 x8.V2.n6 6.93383
R13192 x8.V2.n41 x8.V2.n6 6.93383
R13193 x8.V2.n41 x8.V2.n40 6.93383
R13194 x8.V2.n40 x8.V2.n39 6.93383
R13195 x8.V2.n39 x8.V2.n8 6.93383
R13196 x8.V2.n35 x8.V2.n8 6.93383
R13197 x8.V2.n35 x8.V2.n34 6.93383
R13198 x8.V2.n34 x8.V2.n33 6.93383
R13199 x8.V2.n33 x8.V2.n10 6.93383
R13200 x8.V2.n29 x8.V2.n10 6.93383
R13201 x8.V2.n29 x8.V2.n28 6.93383
R13202 x8.V2.n28 x8.V2.n27 6.93383
R13203 x8.V2.n27 x8.V2.n12 6.93383
R13204 x8.V2.n23 x8.V2.n12 6.93383
R13205 x8.V2.n23 x8.V2.n22 6.93383
R13206 x8.V2.n22 x8.V2.n21 6.93383
R13207 x8.V2.n21 x8.V2.n14 6.93383
R13208 x8.V2.n16 x8.V2.n15 6.93383
R13209 x8.V2.n17 x8.V2.n16 6.93383
R13210 x8.V2.n18 x8.V2.n17 6.93383
R13211 x8.V2.n130 x8.V2.n129 6.86982
R13212 x8.V2.n126 x8.V2.n1 6.47346
R13213 x8.V2.n126 x8.V2.n125 6.27518
R13214 x8.V2.n129 x8.V2.n128 6.23929
R13215 x8.V2.n123 x8.V2.n1 5.09996
R13216 x8.V2.n125 x8.V2.n123 4.87014
R13217 x8.V2.n128 x8.V2.t30 4.35292
R13218 x8.V2.n123 x8.V2.n122 2.7606
R13219 x8.V2.n127 x8.V2 2.58592
R13220 x8.V2.n124 x8.V2.t34 1.45813
R13221 x8.V2.n124 x8.V2.t46 1.45813
R13222 x8.V2.n0 x8.V2.t45 1.45813
R13223 x8.V2.n0 x8.V2.t35 1.45813
R13224 x8.V2.n21 x8.V2.n20 0.7755
R13225 x8.V2.n22 x8.V2.n13 0.7755
R13226 x8.V2.n25 x8.V2.n12 0.7755
R13227 x8.V2.n27 x8.V2.n26 0.7755
R13228 x8.V2.n28 x8.V2.n11 0.7755
R13229 x8.V2.n30 x8.V2.n29 0.7755
R13230 x8.V2.n31 x8.V2.n10 0.7755
R13231 x8.V2.n33 x8.V2.n32 0.7755
R13232 x8.V2.n34 x8.V2.n9 0.7755
R13233 x8.V2.n36 x8.V2.n35 0.7755
R13234 x8.V2.n37 x8.V2.n8 0.7755
R13235 x8.V2.n39 x8.V2.n38 0.7755
R13236 x8.V2.n40 x8.V2.n7 0.7755
R13237 x8.V2.n42 x8.V2.n41 0.7755
R13238 x8.V2.n43 x8.V2.n6 0.7755
R13239 x8.V2.n45 x8.V2.n44 0.7755
R13240 x8.V2.n46 x8.V2.n5 0.7755
R13241 x8.V2.n48 x8.V2.n47 0.7755
R13242 x8.V2.n49 x8.V2.n4 0.7755
R13243 x8.V2.n51 x8.V2.n50 0.7755
R13244 x8.V2.n52 x8.V2.n2 0.7755
R13245 x8.V2.n121 x8.V2.n120 0.7755
R13246 x8.V2.n119 x8.V2.n3 0.7755
R13247 x8.V2.n118 x8.V2.n117 0.7755
R13248 x8.V2.n116 x8.V2.n53 0.7755
R13249 x8.V2.n115 x8.V2.n114 0.7755
R13250 x8.V2.n113 x8.V2.n54 0.7755
R13251 x8.V2.n112 x8.V2.n111 0.7755
R13252 x8.V2.n110 x8.V2.n55 0.7755
R13253 x8.V2.n109 x8.V2.n108 0.7755
R13254 x8.V2.n107 x8.V2.n56 0.7755
R13255 x8.V2.n106 x8.V2.n105 0.7755
R13256 x8.V2.n104 x8.V2.n57 0.7755
R13257 x8.V2.n103 x8.V2.n102 0.7755
R13258 x8.V2.n101 x8.V2.n58 0.7755
R13259 x8.V2.n100 x8.V2.n99 0.7755
R13260 x8.V2.n98 x8.V2.n59 0.7755
R13261 x8.V2.n97 x8.V2.n96 0.7755
R13262 x8.V2.n95 x8.V2.n60 0.7755
R13263 x8.V2.n94 x8.V2.n93 0.7755
R13264 x8.V2.n92 x8.V2.n61 0.7755
R13265 x8.V2.n91 x8.V2.n90 0.7755
R13266 x8.V2.n89 x8.V2.n62 0.7755
R13267 x8.V2.n88 x8.V2.n87 0.7755
R13268 x8.V2.n86 x8.V2.n63 0.7755
R13269 x8.V2.n85 x8.V2.n84 0.7755
R13270 x8.V2.n83 x8.V2.n64 0.7755
R13271 x8.V2.n82 x8.V2.n81 0.7755
R13272 x8.V2.n80 x8.V2.n65 0.7755
R13273 x8.V2.n79 x8.V2.n78 0.7755
R13274 x8.V2.n77 x8.V2.n66 0.7755
R13275 x8.V2.n76 x8.V2.n75 0.7755
R13276 x8.V2.n74 x8.V2.n67 0.7755
R13277 x8.V2.n73 x8.V2.n72 0.7755
R13278 x8.V2.n71 x8.V2.n68 0.7755
R13279 x8.V2.n24 x8.V2.n23 0.7755
R13280 x8.V2.n15 x8.V2.t33 0.763824
R13281 x8.V2.n16 x8.V2.t59 0.763824
R13282 x8.V2.n17 x8.V2.t31 0.763824
R13283 x8.V2.n23 x8.V2.t0 0.763824
R13284 x8.V2.n19 x8.V2.n18 0.684283
R13285 x8.V2.n19 x8.V2.n14 0.629383
R13286 x8.V2.n70 x8.V2.n69 0.629383
R13287 x8.V2 x8.V2.n130 0.403625
R13288 x8.V2.n127 x8.V2.n126 0.219746
R13289 x8.V2.n20 x8.V2.n19 0.145085
R13290 x8.V2.n69 x8.V2.n68 0.145085
R13291 x8.V2.n129 x8.V2.n127 0.0892897
R13292 x8.V2.n20 x8.V2.n13 0.0682083
R13293 x8.V2.n24 x8.V2.n13 0.0682083
R13294 x8.V2.n25 x8.V2.n24 0.0682083
R13295 x8.V2.n26 x8.V2.n25 0.0682083
R13296 x8.V2.n26 x8.V2.n11 0.0682083
R13297 x8.V2.n30 x8.V2.n11 0.0682083
R13298 x8.V2.n31 x8.V2.n30 0.0682083
R13299 x8.V2.n32 x8.V2.n31 0.0682083
R13300 x8.V2.n32 x8.V2.n9 0.0682083
R13301 x8.V2.n36 x8.V2.n9 0.0682083
R13302 x8.V2.n37 x8.V2.n36 0.0682083
R13303 x8.V2.n38 x8.V2.n37 0.0682083
R13304 x8.V2.n38 x8.V2.n7 0.0682083
R13305 x8.V2.n42 x8.V2.n7 0.0682083
R13306 x8.V2.n43 x8.V2.n42 0.0682083
R13307 x8.V2.n44 x8.V2.n43 0.0682083
R13308 x8.V2.n44 x8.V2.n5 0.0682083
R13309 x8.V2.n48 x8.V2.n5 0.0682083
R13310 x8.V2.n49 x8.V2.n48 0.0682083
R13311 x8.V2.n50 x8.V2.n49 0.0682083
R13312 x8.V2.n50 x8.V2.n2 0.0682083
R13313 x8.V2.n121 x8.V2.n3 0.0682083
R13314 x8.V2.n117 x8.V2.n3 0.0682083
R13315 x8.V2.n117 x8.V2.n116 0.0682083
R13316 x8.V2.n116 x8.V2.n115 0.0682083
R13317 x8.V2.n115 x8.V2.n54 0.0682083
R13318 x8.V2.n111 x8.V2.n54 0.0682083
R13319 x8.V2.n111 x8.V2.n110 0.0682083
R13320 x8.V2.n110 x8.V2.n109 0.0682083
R13321 x8.V2.n109 x8.V2.n56 0.0682083
R13322 x8.V2.n105 x8.V2.n56 0.0682083
R13323 x8.V2.n105 x8.V2.n104 0.0682083
R13324 x8.V2.n104 x8.V2.n103 0.0682083
R13325 x8.V2.n103 x8.V2.n58 0.0682083
R13326 x8.V2.n99 x8.V2.n58 0.0682083
R13327 x8.V2.n99 x8.V2.n98 0.0682083
R13328 x8.V2.n98 x8.V2.n97 0.0682083
R13329 x8.V2.n97 x8.V2.n60 0.0682083
R13330 x8.V2.n93 x8.V2.n60 0.0682083
R13331 x8.V2.n93 x8.V2.n92 0.0682083
R13332 x8.V2.n92 x8.V2.n91 0.0682083
R13333 x8.V2.n91 x8.V2.n62 0.0682083
R13334 x8.V2.n87 x8.V2.n62 0.0682083
R13335 x8.V2.n87 x8.V2.n86 0.0682083
R13336 x8.V2.n86 x8.V2.n85 0.0682083
R13337 x8.V2.n85 x8.V2.n64 0.0682083
R13338 x8.V2.n81 x8.V2.n64 0.0682083
R13339 x8.V2.n81 x8.V2.n80 0.0682083
R13340 x8.V2.n80 x8.V2.n79 0.0682083
R13341 x8.V2.n79 x8.V2.n66 0.0682083
R13342 x8.V2.n75 x8.V2.n66 0.0682083
R13343 x8.V2.n75 x8.V2.n74 0.0682083
R13344 x8.V2.n74 x8.V2.n73 0.0682083
R13345 x8.V2.n73 x8.V2.n68 0.0682083
R13346 x8.V2.n122 x8.V2.n121 0.0430347
R13347 x8.V2.n122 x8.V2.n2 0.0256736
R13348 a_12405_n4916.n1 a_12405_n4916.t6 24.0657
R13349 a_12405_n4916.n5 a_12405_n4916.t7 21.5736
R13350 a_12405_n4916.n4 a_12405_n4916.t2 21.5736
R13351 a_12405_n4916.n3 a_12405_n4916.t1 21.5736
R13352 a_12405_n4916.n1 a_12405_n4916.n0 19.6936
R13353 a_12405_n4916.n2 a_12405_n4916.t3 18.5015
R13354 a_12405_n4916.n2 a_12405_n4916.n1 5.46945
R13355 a_12405_n4916.n0 a_12405_n4916.t4 3.55534
R13356 a_12405_n4916.n0 a_12405_n4916.t5 3.55534
R13357 a_12405_n4916.t0 a_12405_n4916.n5 1.60814
R13358 a_12405_n4916.n3 a_12405_n4916.n2 1.04507
R13359 a_12405_n4916.n4 a_12405_n4916.n3 0.0698128
R13360 a_12405_n4916.n5 a_12405_n4916.n4 0.0698128
R13361 a_230_281.t0 a_230_281.t1 37.1785
R13362 a_16157_764.t2 a_16157_764.t0 932.91
R13363 a_16157_764.n6 a_16157_764.t0 361.5
R13364 a_16157_764.n5 a_16157_764.t2 361.5
R13365 a_16157_764.n4 a_16157_764.t6 217.101
R13366 a_16157_764.n4 a_16157_764.t5 216.972
R13367 a_16157_764.n6 a_16157_764.n5 192.569
R13368 a_16157_764.n0 a_16157_764.n4 114.334
R13369 a_16157_764.n5 a_16157_764.n2 80.6505
R13370 a_16157_764.n3 a_16157_764.t4 17.9388
R13371 a_16157_764.n7 a_16157_764.n3 13.5228
R13372 a_16157_764.n3 a_16157_764.n0 2.74902
R13373 a_16157_764.n3 a_16157_764.n2 2.71578
R13374 a_16157_764.t3 a_16157_764.n7 1.84683
R13375 a_16157_764.n7 a_16157_764.t1 1.84683
R13376 a_16157_764.n0 a_16157_764.n1 0.780816
R13377 a_16157_764.n2 a_16157_764.n1 0.165327
R13378 a_16157_764.n6 a_16157_764.n1 80.8153
R13379 a_6605_764.t0 a_6605_764.t2 932.91
R13380 a_6605_764.n6 a_6605_764.t2 361.5
R13381 a_6605_764.n5 a_6605_764.t0 361.5
R13382 a_6605_764.n4 a_6605_764.t5 217.101
R13383 a_6605_764.n4 a_6605_764.t6 216.972
R13384 a_6605_764.n6 a_6605_764.n5 192.569
R13385 a_6605_764.n0 a_6605_764.n4 114.334
R13386 a_6605_764.n5 a_6605_764.n2 80.6505
R13387 a_6605_764.n3 a_6605_764.t4 17.9388
R13388 a_6605_764.n7 a_6605_764.n3 13.5228
R13389 a_6605_764.n3 a_6605_764.n0 2.74902
R13390 a_6605_764.n3 a_6605_764.n2 2.71578
R13391 a_6605_764.n7 a_6605_764.t1 1.84683
R13392 a_6605_764.t3 a_6605_764.n7 1.84683
R13393 a_6605_764.n0 a_6605_764.n1 0.780816
R13394 a_6605_764.n2 a_6605_764.n1 0.165327
R13395 a_6605_764.n6 a_6605_764.n1 80.8153
R13396 a_13817_n9984.n1 a_13817_n9984.t6 24.2695
R13397 a_13817_n9984.n13 a_13817_n9984.t4 21.5736
R13398 a_13817_n9984.n12 a_13817_n9984.t8 21.5736
R13399 a_13817_n9984.n11 a_13817_n9984.t2 21.5736
R13400 a_13817_n9984.n10 a_13817_n9984.t14 21.5736
R13401 a_13817_n9984.n9 a_13817_n9984.t3 21.5736
R13402 a_13817_n9984.n8 a_13817_n9984.t1 21.5736
R13403 a_13817_n9984.n7 a_13817_n9984.t15 21.5736
R13404 a_13817_n9984.n1 a_13817_n9984.n0 19.6768
R13405 a_13817_n9984.n3 a_13817_n9984.n2 19.6768
R13406 a_13817_n9984.n5 a_13817_n9984.n4 19.6768
R13407 a_13817_n9984.n6 a_13817_n9984.t12 18.7802
R13408 a_13817_n9984.n6 a_13817_n9984.n5 5.44609
R13409 a_13817_n9984.n0 a_13817_n9984.t11 3.77447
R13410 a_13817_n9984.n0 a_13817_n9984.t9 3.77447
R13411 a_13817_n9984.n2 a_13817_n9984.t5 3.77447
R13412 a_13817_n9984.n2 a_13817_n9984.t7 3.77447
R13413 a_13817_n9984.n4 a_13817_n9984.t10 3.77447
R13414 a_13817_n9984.n4 a_13817_n9984.t13 3.77447
R13415 a_13817_n9984.t0 a_13817_n9984.n13 1.60814
R13416 a_13817_n9984.n7 a_13817_n9984.n6 1.07925
R13417 a_13817_n9984.n5 a_13817_n9984.n3 0.808313
R13418 a_13817_n9984.n3 a_13817_n9984.n1 0.808313
R13419 a_13817_n9984.n8 a_13817_n9984.n7 0.0698128
R13420 a_13817_n9984.n9 a_13817_n9984.n8 0.0698128
R13421 a_13817_n9984.n10 a_13817_n9984.n9 0.0698128
R13422 a_13817_n9984.n11 a_13817_n9984.n10 0.0698128
R13423 a_13817_n9984.n12 a_13817_n9984.n11 0.0698128
R13424 a_13817_n9984.n13 a_13817_n9984.n12 0.0698128
R13425 a_13817_n4916.n1 a_13817_n4916.t10 24.2695
R13426 a_13817_n4916.n13 a_13817_n4916.t15 21.5736
R13427 a_13817_n4916.n12 a_13817_n4916.t6 21.5736
R13428 a_13817_n4916.n11 a_13817_n4916.t3 21.5736
R13429 a_13817_n4916.n10 a_13817_n4916.t14 21.5736
R13430 a_13817_n4916.n9 a_13817_n4916.t1 21.5736
R13431 a_13817_n4916.n8 a_13817_n4916.t4 21.5736
R13432 a_13817_n4916.n7 a_13817_n4916.t2 21.5736
R13433 a_13817_n4916.n1 a_13817_n4916.n0 19.6768
R13434 a_13817_n4916.n3 a_13817_n4916.n2 19.6768
R13435 a_13817_n4916.n5 a_13817_n4916.n4 19.6768
R13436 a_13817_n4916.n6 a_13817_n4916.t11 18.7802
R13437 a_13817_n4916.n6 a_13817_n4916.n5 5.44609
R13438 a_13817_n4916.n0 a_13817_n4916.t7 3.77447
R13439 a_13817_n4916.n0 a_13817_n4916.t8 3.77447
R13440 a_13817_n4916.n2 a_13817_n4916.t5 3.77447
R13441 a_13817_n4916.n2 a_13817_n4916.t12 3.77447
R13442 a_13817_n4916.n4 a_13817_n4916.t9 3.77447
R13443 a_13817_n4916.n4 a_13817_n4916.t13 3.77447
R13444 a_13817_n4916.t0 a_13817_n4916.n13 1.60814
R13445 a_13817_n4916.n7 a_13817_n4916.n6 1.07925
R13446 a_13817_n4916.n5 a_13817_n4916.n3 0.808313
R13447 a_13817_n4916.n3 a_13817_n4916.n1 0.808313
R13448 a_13817_n4916.n8 a_13817_n4916.n7 0.0698128
R13449 a_13817_n4916.n9 a_13817_n4916.n8 0.0698128
R13450 a_13817_n4916.n10 a_13817_n4916.n9 0.0698128
R13451 a_13817_n4916.n11 a_13817_n4916.n10 0.0698128
R13452 a_13817_n4916.n12 a_13817_n4916.n11 0.0698128
R13453 a_13817_n4916.n13 a_13817_n4916.n12 0.0698128
R13454 D9.n3 D9.t2 186.374
R13455 D9.n2 D9.n1 184.464
R13456 D9.n3 D9.t1 170.308
R13457 D9.n4 D9.n3 165.827
R13458 D9.n0 D9.t0 46.372
R13459 D9.n4 D9.n2 13.2781
R13460 D9.n2 D9 5.71063
R13461 D9.n1 D9 4.3525
R13462 D9 D9.n0 3.61505
R13463 D9.n0 D9 2.5677
R13464 D9.n1 D9 1.96317
R13465 D9 D9.n4 1.24229
R13466 D63v3.n4 D63v3.n3 873.303
R13467 D63v3 D63v3.n4 585
R13468 D63v3.t1 D63v3 506.99
R13469 D63v3 D63v3.t0 150.315
R13470 D63v3.n4 D63v3.t1 147.756
R13471 D63v3.n1 D63v3.t3 110.788
R13472 D63v3.n0 D63v3.t2 110.698
R13473 D63v3.n0 D63v3.t4 110.397
R13474 D63v3.n2 D63v3.t5 105.519
R13475 D63v3 D63v3.n0 22.9067
R13476 D63v3.n0 D63v3.n2 8.99346
R13477 D63v3.n1 D63v3 7.10988
R13478 D63v3.n0 D63v3 6.99737
R13479 D63v3.n3 D63v3 4.99562
R13480 D63v3.n2 D63v3.n1 4.88025
R13481 D63v3 D63v3.n3 2.70619
R13482 a_16150_281.t0 a_16150_281.t1 37.1785
R13483 a_12973_764.t0 a_12973_764.t2 932.91
R13484 a_12973_764.n6 a_12973_764.t2 361.5
R13485 a_12973_764.n5 a_12973_764.t0 361.5
R13486 a_12973_764.n4 a_12973_764.t5 217.101
R13487 a_12973_764.n4 a_12973_764.t6 216.972
R13488 a_12973_764.n6 a_12973_764.n5 192.569
R13489 a_12973_764.n0 a_12973_764.n4 114.334
R13490 a_12973_764.n5 a_12973_764.n2 80.6505
R13491 a_12973_764.n3 a_12973_764.t4 17.9388
R13492 a_12973_764.n7 a_12973_764.n3 13.5228
R13493 a_12973_764.n3 a_12973_764.n0 2.74902
R13494 a_12973_764.n3 a_12973_764.n2 2.71578
R13495 a_12973_764.n7 a_12973_764.t1 1.84683
R13496 a_12973_764.t3 a_12973_764.n7 1.84683
R13497 a_12973_764.n0 a_12973_764.n1 0.780816
R13498 a_12973_764.n2 a_12973_764.n1 0.165327
R13499 a_12973_764.n6 a_12973_764.n1 80.8153
R13500 D03v3.n3 D03v3.n2 873.303
R13501 D03v3 D03v3.n3 585
R13502 D03v3.t1 D03v3 506.99
R13503 D03v3 D03v3.t0 150.315
R13504 D03v3.n3 D03v3.t1 147.756
R13505 D03v3.n0 D03v3.t2 104.644
R13506 D03v3.n1 D03v3.t3 104.257
R13507 D03v3.n1 D03v3.n0 13.3986
R13508 D03v3.n0 D03v3 10.6402
R13509 D03v3 D03v3.n1 6.12044
R13510 D03v3.n2 D03v3 4.99562
R13511 D03v3 D03v3.n2 2.70619
R13512 a_10583_764.t5 a_10583_764.n1 553.975
R13513 a_10583_764.n6 a_10583_764.t5 553.975
R13514 a_10583_764.n5 a_10583_764.t6 275.969
R13515 a_10583_764.n3 a_10583_764.t4 275.969
R13516 a_10583_764.n4 a_10583_764.t7 275.877
R13517 a_10583_764.n9 a_10583_764.t3 15.8632
R13518 a_10583_764.n10 a_10583_764.n9 13.5228
R13519 a_10583_764.n9 a_10583_764.n8 5.588
R13520 a_10583_764.n7 a_10583_764.n6 2.79633
R13521 a_10583_764.n8 a_10583_764.n7 2.52001
R13522 a_10583_764.n3 a_10583_764.n0 2.34014
R13523 a_10583_764.n2 a_10583_764.n3 2.3327
R13524 a_10583_764.n2 a_10583_764.n4 2.23523
R13525 a_10583_764.n4 a_10583_764.n0 2.23295
R13526 a_10583_764.n5 a_10583_764.n2 2.04972
R13527 a_10583_764.n0 a_10583_764.n5 2.04764
R13528 a_10583_764.t0 a_10583_764.n10 1.84683
R13529 a_10583_764.n10 a_10583_764.t1 1.84683
R13530 a_10583_764.n8 a_10583_764.t2 1.73283
R13531 a_10583_764.n7 a_10583_764.n1 1.29633
R13532 a_10583_764.n6 a_10583_764.n0 0.585777
R13533 a_10583_764.n2 a_10583_764.n1 0.569287
R13534 a_204_12823.n3 a_204_12823.t9 230.883
R13535 a_204_12823.n0 a_204_12823.t6 230.883
R13536 a_204_12823.n3 a_204_12823.t8 230.363
R13537 a_204_12823.n3 a_204_12823.t7 230.363
R13538 a_204_12823.n4 a_204_12823.t5 230.363
R13539 a_204_12823.n4 a_204_12823.t12 230.363
R13540 a_204_12823.n2 a_204_12823.t11 230.363
R13541 a_204_12823.n2 a_204_12823.t10 230.363
R13542 a_204_12823.n2 a_204_12823.t14 230.363
R13543 a_204_12823.n1 a_204_12823.t13 230.363
R13544 a_204_12823.n1 a_204_12823.t16 230.363
R13545 a_204_12823.n0 a_204_12823.t15 230.363
R13546 a_204_12823.n6 a_204_12823.t4 227.346
R13547 a_204_12823.n7 a_204_12823.t2 227.346
R13548 a_204_12823.n5 a_204_12823.t1 60.2247
R13549 a_204_12823.n5 a_204_12823.t3 60.2247
R13550 a_204_12823.t0 a_204_12823.n8 7.89252
R13551 a_204_12823.n5 a_204_12823.n2 4.10301
R13552 a_204_12823.n8 a_204_12823.n7 2.88104
R13553 a_204_12823.n8 a_204_12823.n6 2.49107
R13554 a_204_12823.n2 a_204_12823.n4 1.56098
R13555 a_204_12823.n5 a_204_12823.n6 1.33032
R13556 a_204_12823.n7 a_204_12823.n5 1.11879
R13557 a_204_12823.n4 a_204_12823.n3 1.04082
R13558 a_204_12823.n2 a_204_12823.n1 1.04082
R13559 a_204_12823.n1 a_204_12823.n0 1.04082
R13560 a_9789_764.t1 a_9789_764.t3 932.91
R13561 a_9789_764.n6 a_9789_764.t3 361.5
R13562 a_9789_764.n5 a_9789_764.t1 361.5
R13563 a_9789_764.n2 a_9789_764.t5 217.101
R13564 a_9789_764.n2 a_9789_764.t6 216.972
R13565 a_9789_764.n6 a_9789_764.n5 192.569
R13566 a_9789_764.n3 a_9789_764.n2 114.334
R13567 a_9789_764.n7 a_9789_764.n6 80.6505
R13568 a_9789_764.n5 a_9789_764.n4 80.6505
R13569 a_9789_764.n0 a_9789_764.t0 17.9388
R13570 a_9789_764.n9 a_9789_764.n0 13.5228
R13571 a_9789_764.n0 a_9789_764.n8 2.74902
R13572 a_9789_764.n0 a_9789_764.n1 2.71578
R13573 a_9789_764.n9 a_9789_764.t2 1.84683
R13574 a_9789_764.t4 a_9789_764.n9 1.84683
R13575 a_9789_764.n8 a_9789_764.n7 1.72446
R13576 a_9789_764.n4 a_9789_764.n3 1.5005
R13577 a_9789_764.n8 a_9789_764.n3 0.224458
R13578 a_9789_764.n7 a_9789_764.n1 0.182141
R13579 a_9789_764.n4 a_9789_764.n1 0.182141
R13580 ia_opamp_0.ibias.n6 ia_opamp_0.ibias.t5 281.942
R13581 ia_opamp_0.ibias.n3 ia_opamp_0.ibias.t4 232.155
R13582 ia_opamp_0.ibias.n4 ia_opamp_0.ibias.t0 232.155
R13583 ia_opamp_0.ibias ia_opamp_0.ibias.n2 15.9991
R13584 ia_opamp_0.ibias ia_opamp_0.ibias.n1 15.4767
R13585 ia_opamp_0.ibias.n5 ia_opamp_0.ibias.t1 5.4926
R13586 ia_opamp_0.ibias.n0 ia_opamp_0.ibias.n3 4.11682
R13587 ia_opamp_0.ibias.n3 ia_opamp_0.ibias.n1 4.11576
R13588 ia_opamp_0.ibias.n0 ia_opamp_0.ibias.n4 3.20309
R13589 ia_opamp_0.ibias.n4 ia_opamp_0.ibias.n1 3.20309
R13590 ia_opamp_0.ibias.n5 ia_opamp_0.ibias.n0 2.71404
R13591 ia_opamp_0.ibias.n2 ia_opamp_0.ibias.t3 1.84683
R13592 ia_opamp_0.ibias.n2 ia_opamp_0.ibias.t2 1.84683
R13593 ia_opamp_0.ibias.n6 ia_opamp_0.ibias.n5 1.5165
R13594 ia_opamp_0.ibias.n1 ia_opamp_0.ibias.n6 0.960738
R13595 ia_opamp_0.ibias.n0 ia_opamp_0.ibias 0.953625
R13596 D3.n3 D3.t2 186.374
R13597 D3.n2 D3.n1 184.464
R13598 D3.n3 D3.t0 170.308
R13599 D3.n4 D3.n3 165.827
R13600 D3.n0 D3.t1 46.372
R13601 D3.n4 D3.n2 13.2781
R13602 D3.n2 D3 5.71063
R13603 D3.n1 D3 4.3525
R13604 D3 D3.n0 3.61505
R13605 D3.n0 D3 2.5677
R13606 D3.n1 D3 1.96317
R13607 D3 D3.n4 1.24229
R13608 D5.n3 D5.t2 186.374
R13609 D5.n2 D5.n1 184.464
R13610 D5.n3 D5.t0 170.308
R13611 D5.n4 D5.n3 165.827
R13612 D5.n0 D5.t1 46.372
R13613 D5.n4 D5.n2 13.2781
R13614 D5.n2 D5 5.71063
R13615 D5.n1 D5 4.3525
R13616 D5 D5.n0 3.61505
R13617 D5.n0 D5 2.5677
R13618 D5.n1 D5 1.96317
R13619 D5 D5.n4 1.24229
R13620 D4.n3 D4.t2 186.374
R13621 D4.n2 D4.n1 184.464
R13622 D4.n3 D4.t0 170.308
R13623 D4.n4 D4.n3 165.827
R13624 D4.n0 D4.t1 46.372
R13625 D4.n4 D4.n2 13.2781
R13626 D4.n2 D4 5.71063
R13627 D4.n1 D4 4.3525
R13628 D4 D4.n0 3.61505
R13629 D4.n0 D4 2.5677
R13630 D4.n1 D4 1.96317
R13631 D4 D4.n4 1.24229
R13632 amp_biases_0.ibias1.n7 amp_biases_0.ibias1.t4 281.421
R13633 amp_biases_0.ibias1.n3 amp_biases_0.ibias1.t5 232.155
R13634 amp_biases_0.ibias1.n4 amp_biases_0.ibias1.t0 232.155
R13635 amp_biases_0.ibias1 amp_biases_0.ibias1.n7 20.3794
R13636 amp_biases_0.ibias1 amp_biases_0.ibias1.n1 15.9991
R13637 amp_biases_0.ibias1.n5 amp_biases_0.ibias1.t1 5.4926
R13638 amp_biases_0.ibias1.n0 amp_biases_0.ibias1.n3 4.11682
R13639 amp_biases_0.ibias1.n3 amp_biases_0.ibias1.n2 4.11576
R13640 amp_biases_0.ibias1.n4 amp_biases_0.ibias1.n2 3.20309
R13641 amp_biases_0.ibias1.n0 amp_biases_0.ibias1.n4 3.20309
R13642 amp_biases_0.ibias1.n5 amp_biases_0.ibias1.n0 2.71404
R13643 amp_biases_0.ibias1.n1 amp_biases_0.ibias1.t3 1.84683
R13644 amp_biases_0.ibias1.n1 amp_biases_0.ibias1.t2 1.84683
R13645 amp_biases_0.ibias1.n6 amp_biases_0.ibias1.n5 1.50744
R13646 amp_biases_0.ibias1.n6 amp_biases_0.ibias1.n2 1.19321
R13647 amp_biases_0.ibias1.n0 amp_biases_0.ibias1 0.953625
R13648 amp_biases_0.ibias1.n7 amp_biases_0.ibias1.n6 0.531297
R13649 a_10047_764.n0 a_10047_764.t1 6.15493
R13650 a_10047_764.n0 a_10047_764.t2 5.15685
R13651 a_10047_764.t0 a_10047_764.n0 5.15662
R13652 a_3421_764.t3 a_3421_764.t1 932.91
R13653 a_3421_764.n6 a_3421_764.t1 361.5
R13654 a_3421_764.n5 a_3421_764.t3 361.5
R13655 a_3421_764.n4 a_3421_764.t6 217.101
R13656 a_3421_764.n4 a_3421_764.t5 216.972
R13657 a_3421_764.n6 a_3421_764.n5 192.569
R13658 a_3421_764.n0 a_3421_764.n4 114.334
R13659 a_3421_764.n5 a_3421_764.n2 80.6505
R13660 a_3421_764.n3 a_3421_764.t0 17.9388
R13661 a_3421_764.n7 a_3421_764.n3 13.5228
R13662 a_3421_764.n3 a_3421_764.n0 2.74902
R13663 a_3421_764.n3 a_3421_764.n2 2.71578
R13664 a_3421_764.t4 a_3421_764.n7 1.84683
R13665 a_3421_764.n7 a_3421_764.t2 1.84683
R13666 a_3421_764.n0 a_3421_764.n1 0.780816
R13667 a_3421_764.n2 a_3421_764.n1 0.165327
R13668 a_3421_764.n6 a_3421_764.n1 80.8153
R13669 a_4215_764.t7 a_4215_764.n0 553.975
R13670 a_4215_764.n8 a_4215_764.t7 553.975
R13671 a_4215_764.n6 a_4215_764.t6 275.969
R13672 a_4215_764.n2 a_4215_764.t4 275.969
R13673 a_4215_764.n3 a_4215_764.t5 275.877
R13674 a_4215_764.n11 a_4215_764.t0 15.8632
R13675 a_4215_764.n12 a_4215_764.n11 13.5228
R13676 a_4215_764.n11 a_4215_764.n10 5.588
R13677 a_4215_764.n9 a_4215_764.n8 2.79633
R13678 a_4215_764.n10 a_4215_764.n9 2.52001
R13679 a_4215_764.n2 a_4215_764.n1 2.34014
R13680 a_4215_764.n4 a_4215_764.n2 2.3327
R13681 a_4215_764.n4 a_4215_764.n3 2.23523
R13682 a_4215_764.n3 a_4215_764.n1 2.23295
R13683 a_4215_764.n6 a_4215_764.n5 2.04972
R13684 a_4215_764.n7 a_4215_764.n6 2.04764
R13685 a_4215_764.n12 a_4215_764.t2 1.84683
R13686 a_4215_764.t3 a_4215_764.n12 1.84683
R13687 a_4215_764.n10 a_4215_764.t1 1.73283
R13688 a_4215_764.n9 a_4215_764.n0 1.29633
R13689 a_4215_764.n8 a_4215_764.n7 0.295289
R13690 a_4215_764.n7 a_4215_764.n1 0.290988
R13691 a_4215_764.n5 a_4215_764.n0 0.288208
R13692 a_4215_764.n5 a_4215_764.n4 0.281579
R13693 a_237_764.t2 a_237_764.t0 932.91
R13694 a_237_764.n6 a_237_764.t0 361.5
R13695 a_237_764.n5 a_237_764.t2 361.5
R13696 a_237_764.n4 a_237_764.t5 217.101
R13697 a_237_764.n4 a_237_764.t6 216.972
R13698 a_237_764.n6 a_237_764.n5 192.569
R13699 a_237_764.n0 a_237_764.n4 114.334
R13700 a_237_764.n5 a_237_764.n2 80.6505
R13701 a_237_764.n3 a_237_764.t4 17.9388
R13702 a_237_764.n7 a_237_764.n3 13.5228
R13703 a_237_764.n3 a_237_764.n0 2.74902
R13704 a_237_764.n3 a_237_764.n2 2.71578
R13705 a_237_764.t3 a_237_764.n7 1.84683
R13706 a_237_764.n7 a_237_764.t1 1.84683
R13707 a_237_764.n0 a_237_764.n1 0.780816
R13708 a_237_764.n2 a_237_764.n1 0.165327
R13709 a_237_764.n6 a_237_764.n1 80.8153
R13710 a_495_764.n0 a_495_764.t1 6.15493
R13711 a_495_764.t0 a_495_764.n0 5.15685
R13712 a_495_764.n0 a_495_764.t2 5.15662
R13713 a_7399_764.t5 a_7399_764.n0 553.975
R13714 a_7399_764.n8 a_7399_764.t5 553.975
R13715 a_7399_764.n6 a_7399_764.t7 275.969
R13716 a_7399_764.n2 a_7399_764.t4 275.969
R13717 a_7399_764.n3 a_7399_764.t6 275.877
R13718 a_7399_764.n11 a_7399_764.t3 15.8632
R13719 a_7399_764.n12 a_7399_764.n11 13.5228
R13720 a_7399_764.n11 a_7399_764.n10 5.588
R13721 a_7399_764.n9 a_7399_764.n8 2.79633
R13722 a_7399_764.n10 a_7399_764.n9 2.52001
R13723 a_7399_764.n2 a_7399_764.n1 2.34014
R13724 a_7399_764.n4 a_7399_764.n2 2.3327
R13725 a_7399_764.n4 a_7399_764.n3 2.23523
R13726 a_7399_764.n3 a_7399_764.n1 2.23295
R13727 a_7399_764.n6 a_7399_764.n5 2.04972
R13728 a_7399_764.n7 a_7399_764.n6 2.04764
R13729 a_7399_764.t1 a_7399_764.n12 1.84683
R13730 a_7399_764.n12 a_7399_764.t0 1.84683
R13731 a_7399_764.n10 a_7399_764.t2 1.73283
R13732 a_7399_764.n9 a_7399_764.n0 1.29633
R13733 a_7399_764.n8 a_7399_764.n7 0.295289
R13734 a_7399_764.n7 a_7399_764.n1 0.290988
R13735 a_7399_764.n5 a_7399_764.n0 0.288208
R13736 a_7399_764.n5 a_7399_764.n4 0.281579
R13737 D2.n3 D2.t2 186.374
R13738 D2.n2 D2.n1 184.464
R13739 D2.n3 D2.t0 170.308
R13740 D2.n4 D2.n3 165.827
R13741 D2.n0 D2.t1 46.372
R13742 D2.n4 D2.n2 13.2781
R13743 D2.n2 D2 5.71063
R13744 D2.n1 D2 4.3525
R13745 D2 D2.n0 3.61505
R13746 D2.n0 D2 2.5677
R13747 D2.n1 D2 1.96317
R13748 D2 D2.n4 1.24229
R13749 V2.n0 V2.t0 492.844
R13750 V2.n0 V2 4.95011
R13751 V2 V2.n0 0.063
R13752 a_3679_764.n0 a_3679_764.t0 6.15493
R13753 a_3679_764.n0 a_3679_764.t2 5.15685
R13754 a_3679_764.t1 a_3679_764.n0 5.15662
R13755 D53v3.n3 D53v3.n2 873.303
R13756 D53v3 D53v3.n3 585
R13757 D53v3.t1 D53v3 506.99
R13758 D53v3 D53v3.t0 150.315
R13759 D53v3.n3 D53v3.t1 147.756
R13760 D53v3.n0 D53v3.t2 109.188
R13761 D53v3.n1 D53v3.t3 104.257
R13762 D53v3 D53v3.n0 21.9036
R13763 D53v3.n1 D53v3 11.0267
R13764 D53v3.n0 D53v3 8.4231
R13765 D53v3.n0 D53v3.n1 6.51308
R13766 D53v3.n2 D53v3 4.99562
R13767 D53v3 D53v3.n2 2.70619
R13768 G.n0 G.t0 492.887
R13769 G.n0 G 6.0151
R13770 G G.n0 0.01925
R13771 D13v3.n5 D13v3.n4 873.303
R13772 D13v3 D13v3.n5 585
R13773 D13v3.t1 D13v3 506.99
R13774 D13v3 D13v3.t0 150.315
R13775 D13v3.n5 D13v3.t1 147.756
R13776 D13v3.n1 D13v3.t2 110.788
R13777 D13v3.n0 D13v3.t3 110.788
R13778 D13v3.n2 D13v3.t4 105.791
R13779 D13v3.n3 D13v3.t5 105.519
R13780 D13v3.n3 D13v3.n2 13.3894
R13781 D13v3.n1 D13v3 7.10988
R13782 D13v3.n4 D13v3 4.99562
R13783 D13v3.n0 D13v3.n3 4.87929
R13784 D13v3.n2 D13v3.n1 4.60644
R13785 D13v3 D13v3.n0 3.39112
R13786 D13v3 D13v3.n4 2.70619
R13787 D7.n3 D7.t2 186.374
R13788 D7.n2 D7.n1 184.464
R13789 D7.n3 D7.t1 170.308
R13790 D7.n4 D7.n3 165.827
R13791 D7.n0 D7.t0 46.372
R13792 D7.n4 D7.n2 13.2781
R13793 D7.n2 D7 5.71063
R13794 D7.n1 D7 4.3525
R13795 D7 D7.n0 3.61505
R13796 D7.n0 D7 2.5677
R13797 D7.n1 D7 1.96317
R13798 D7 D7.n4 1.24229
R13799 amp_biases_0.ibias5.n5 amp_biases_0.ibias5.t4 281.947
R13800 amp_biases_0.ibias5.n2 amp_biases_0.ibias5.t5 232.155
R13801 amp_biases_0.ibias5.n3 amp_biases_0.ibias5.t0 232.155
R13802 amp_biases_0.ibias5 amp_biases_0.ibias5.n1 22.7505
R13803 amp_biases_0.ibias5 amp_biases_0.ibias5.n6 15.9408
R13804 amp_biases_0.ibias5.n4 amp_biases_0.ibias5.t1 5.4926
R13805 amp_biases_0.ibias5.n0 amp_biases_0.ibias5.n2 4.11682
R13806 amp_biases_0.ibias5.n2 amp_biases_0.ibias5.n1 4.11576
R13807 amp_biases_0.ibias5.n0 amp_biases_0.ibias5.n3 3.20309
R13808 amp_biases_0.ibias5.n3 amp_biases_0.ibias5.n1 3.20309
R13809 amp_biases_0.ibias5.n4 amp_biases_0.ibias5.n0 2.71404
R13810 amp_biases_0.ibias5.n6 amp_biases_0.ibias5.t3 1.84683
R13811 amp_biases_0.ibias5.n6 amp_biases_0.ibias5.t2 1.84683
R13812 amp_biases_0.ibias5.n5 amp_biases_0.ibias5.n4 1.51107
R13813 amp_biases_0.ibias5.n1 amp_biases_0.ibias5.n5 1.07882
R13814 amp_biases_0.ibias5.n0 amp_biases_0.ibias5 0.953625
R13815 D23v3.n5 D23v3.n4 873.303
R13816 D23v3 D23v3.n5 585
R13817 D23v3.t1 D23v3 506.99
R13818 D23v3 D23v3.t0 150.315
R13819 D23v3.n5 D23v3.t1 147.756
R13820 D23v3.n1 D23v3.t8 108.13
R13821 D23v3.n0 D23v3.t9 108.13
R13822 D23v3.n1 D23v3.t6 107.737
R13823 D23v3.n1 D23v3.t4 107.737
R13824 D23v3.n0 D23v3.t7 107.737
R13825 D23v3.n0 D23v3.t5 107.737
R13826 D23v3.n2 D23v3.t2 103.1
R13827 D23v3.n3 D23v3.t3 102.909
R13828 D23v3.n3 D23v3.n2 13.4096
R13829 D23v3.n1 D23v3 8.5005
R13830 D23v3 D23v3.n0 5.588
R13831 D23v3.n2 D23v3.n1 5.44346
R13832 D23v3.n4 D23v3 4.99562
R13833 D23v3.n0 D23v3.n3 4.82852
R13834 D23v3 D23v3.n4 2.70619
R13835 a_2308_n9984.n1 a_2308_n9984.t3 24.0657
R13836 a_2308_n9984.n3 a_2308_n9984.t6 21.6429
R13837 a_2308_n9984.n3 a_2308_n9984.t7 21.5736
R13838 a_2308_n9984.n4 a_2308_n9984.t5 21.5736
R13839 a_2308_n9984.n1 a_2308_n9984.n0 19.6936
R13840 a_2308_n9984.n2 a_2308_n9984.t0 18.5015
R13841 a_2308_n9984.n2 a_2308_n9984.n1 5.46945
R13842 a_2308_n9984.n0 a_2308_n9984.t2 3.55534
R13843 a_2308_n9984.n0 a_2308_n9984.t1 3.55534
R13844 a_2308_n9984.t4 a_2308_n9984.n5 1.53882
R13845 a_2308_n9984.n5 a_2308_n9984.n2 1.04507
R13846 a_2308_n9984.n5 a_2308_n9984.n4 0.0698128
R13847 a_2308_n9984.n4 a_2308_n9984.n3 0.0698128
R13848 a_2308_n4916.n1 a_2308_n4916.t3 24.0657
R13849 a_2308_n4916.n3 a_2308_n4916.t6 21.6429
R13850 a_2308_n4916.n3 a_2308_n4916.t5 21.5736
R13851 a_2308_n4916.n4 a_2308_n4916.t7 21.5736
R13852 a_2308_n4916.n1 a_2308_n4916.n0 19.6936
R13853 a_2308_n4916.n2 a_2308_n4916.t0 18.5015
R13854 a_2308_n4916.n2 a_2308_n4916.n1 5.46945
R13855 a_2308_n4916.n0 a_2308_n4916.t2 3.55534
R13856 a_2308_n4916.n0 a_2308_n4916.t1 3.55534
R13857 a_2308_n4916.t4 a_2308_n4916.n5 1.53882
R13858 a_2308_n4916.n5 a_2308_n4916.n2 1.04507
R13859 a_2308_n4916.n5 a_2308_n4916.n4 0.0698128
R13860 a_2308_n4916.n4 a_2308_n4916.n3 0.0698128
R13861 amp_biases_0.ibias2.n6 amp_biases_0.ibias2.t5 281.421
R13862 amp_biases_0.ibias2.n2 amp_biases_0.ibias2.t4 232.155
R13863 amp_biases_0.ibias2.n3 amp_biases_0.ibias2.t0 232.155
R13864 amp_biases_0.ibias2 amp_biases_0.ibias2.n6 21.0783
R13865 amp_biases_0.ibias2 amp_biases_0.ibias2.n7 19.9252
R13866 amp_biases_0.ibias2.n4 amp_biases_0.ibias2.t1 5.4926
R13867 amp_biases_0.ibias2.n0 amp_biases_0.ibias2.n2 4.11682
R13868 amp_biases_0.ibias2.n2 amp_biases_0.ibias2.n1 4.11576
R13869 amp_biases_0.ibias2.n3 amp_biases_0.ibias2.n1 3.20309
R13870 amp_biases_0.ibias2.n0 amp_biases_0.ibias2.n3 3.20309
R13871 amp_biases_0.ibias2.n4 amp_biases_0.ibias2.n0 2.71404
R13872 amp_biases_0.ibias2.n7 amp_biases_0.ibias2.t3 1.84683
R13873 amp_biases_0.ibias2.n7 amp_biases_0.ibias2.t2 1.84683
R13874 amp_biases_0.ibias2.n5 amp_biases_0.ibias2.n4 1.50744
R13875 amp_biases_0.ibias2.n5 amp_biases_0.ibias2.n1 1.19321
R13876 amp_biases_0.ibias2.n0 amp_biases_0.ibias2 0.953625
R13877 amp_biases_0.ibias2.n6 amp_biases_0.ibias2.n5 0.531297
R13878 a_3414_281.t0 a_3414_281.t1 37.1785
R13879 D1.n3 D1.t2 186.374
R13880 D1.n2 D1.n1 184.464
R13881 D1.n3 D1.t0 170.308
R13882 D1.n4 D1.n3 165.827
R13883 D1.n0 D1.t1 46.372
R13884 D1.n4 D1.n2 13.2781
R13885 D1.n2 D1 5.71063
R13886 D1.n1 D1 4.3525
R13887 D1 D1.n0 3.61505
R13888 D1.n0 D1 2.5677
R13889 D1.n1 D1 1.96317
R13890 D1 D1.n4 1.24229
R13891 a_13767_764.t5 a_13767_764.n0 553.975
R13892 a_13767_764.n8 a_13767_764.t5 553.975
R13893 a_13767_764.n6 a_13767_764.t4 275.969
R13894 a_13767_764.n2 a_13767_764.t7 275.969
R13895 a_13767_764.n3 a_13767_764.t6 275.877
R13896 a_13767_764.n11 a_13767_764.t3 15.8632
R13897 a_13767_764.n12 a_13767_764.n11 13.5228
R13898 a_13767_764.n11 a_13767_764.n10 5.588
R13899 a_13767_764.n9 a_13767_764.n8 2.79633
R13900 a_13767_764.n10 a_13767_764.n9 2.52001
R13901 a_13767_764.n2 a_13767_764.n1 2.34014
R13902 a_13767_764.n4 a_13767_764.n2 2.3327
R13903 a_13767_764.n4 a_13767_764.n3 2.23523
R13904 a_13767_764.n3 a_13767_764.n1 2.23295
R13905 a_13767_764.n6 a_13767_764.n5 2.04972
R13906 a_13767_764.n7 a_13767_764.n6 2.04764
R13907 a_13767_764.t1 a_13767_764.n12 1.84683
R13908 a_13767_764.n12 a_13767_764.t0 1.84683
R13909 a_13767_764.n10 a_13767_764.t2 1.73283
R13910 a_13767_764.n9 a_13767_764.n0 1.29633
R13911 a_13767_764.n8 a_13767_764.n7 0.295289
R13912 a_13767_764.n7 a_13767_764.n1 0.290988
R13913 a_13767_764.n5 a_13767_764.n0 0.288208
R13914 a_13767_764.n5 a_13767_764.n4 0.281579
R13915 a_6863_764.n0 a_6863_764.t0 6.15493
R13916 a_6863_764.t1 a_6863_764.n0 5.15685
R13917 a_6863_764.n0 a_6863_764.t2 5.15662
R13918 a_6598_281.t0 a_6598_281.t1 37.1785
R13919 D0.n3 D0.t2 186.374
R13920 D0.n2 D0.n1 184.464
R13921 D0.n3 D0.t0 170.308
R13922 D0.n4 D0.n3 165.827
R13923 D0.n0 D0.t1 46.372
R13924 D0.n4 D0.n2 13.2781
R13925 D0.n2 D0 5.71063
R13926 D0.n1 D0 4.3525
R13927 D0 D0.n0 3.61505
R13928 D0.n0 D0 2.5677
R13929 D0.n1 D0 1.96317
R13930 D0 D0.n4 1.24229
R13931 sky130_fd_sc_hvl__lsbuflv2hv_1_0[10].X.n2 sky130_fd_sc_hvl__lsbuflv2hv_1_0[10].X.n1 873.303
R13932 sky130_fd_sc_hvl__lsbuflv2hv_1_0[10].X sky130_fd_sc_hvl__lsbuflv2hv_1_0[10].X.n2 585
R13933 sky130_fd_sc_hvl__lsbuflv2hv_1_0[10].X.t1 sky130_fd_sc_hvl__lsbuflv2hv_1_0[10].X 506.99
R13934 sky130_fd_sc_hvl__lsbuflv2hv_1_0[10].X.n0 sky130_fd_sc_hvl__lsbuflv2hv_1_0[10].X.t2 235.912
R13935 sky130_fd_sc_hvl__lsbuflv2hv_1_0[10].X.n0 sky130_fd_sc_hvl__lsbuflv2hv_1_0[10].X.t3 235.048
R13936 sky130_fd_sc_hvl__lsbuflv2hv_1_0[10].X sky130_fd_sc_hvl__lsbuflv2hv_1_0[10].X.t0 150.315
R13937 sky130_fd_sc_hvl__lsbuflv2hv_1_0[10].X.n2 sky130_fd_sc_hvl__lsbuflv2hv_1_0[10].X.t1 147.756
R13938 sky130_fd_sc_hvl__lsbuflv2hv_1_0[10].X sky130_fd_sc_hvl__lsbuflv2hv_1_0[10].X.n0 6.98521
R13939 sky130_fd_sc_hvl__lsbuflv2hv_1_0[10].X.n1 sky130_fd_sc_hvl__lsbuflv2hv_1_0[10].X 4.99562
R13940 sky130_fd_sc_hvl__lsbuflv2hv_1_0[10].X sky130_fd_sc_hvl__lsbuflv2hv_1_0[10].X.n1 2.70619
R13941 a_2622_12748.n0 a_2622_12748.t3 235.228
R13942 a_2622_12748.n0 a_2622_12748.t1 234.392
R13943 a_2622_12748.n1 a_2622_12748.n0 7.01736
R13944 a_2622_12748.n1 a_2622_12748.t0 1.0711
R13945 a_2622_12748.t2 a_2622_12748.n1 1.0711
R13946 ibias ibias.t0 8.20856
R13947 a_12966_281.t0 a_12966_281.t1 37.1785
R13948 ena.n3 ena.t2 186.374
R13949 ena.n2 ena.n1 184.464
R13950 ena.n3 ena.t1 170.308
R13951 ena.n4 ena.n3 165.827
R13952 ena.n0 ena.t0 46.372
R13953 ena.n4 ena.n2 13.2781
R13954 ena.n2 ena 5.71063
R13955 ena.n1 ena 4.3525
R13956 ena ena.n0 3.61505
R13957 ena.n0 ena 2.5677
R13958 ena.n1 ena 1.96317
R13959 ena ena.n4 1.24229
R13960 a_9782_281.t0 a_9782_281.t1 37.1785
R13961 amp_biases_0.ibias3.n6 amp_biases_0.ibias3.t5 281.421
R13962 amp_biases_0.ibias3.n2 amp_biases_0.ibias3.t4 232.155
R13963 amp_biases_0.ibias3.n3 amp_biases_0.ibias3.t0 232.155
R13964 amp_biases_0.ibias3 amp_biases_0.ibias3.n6 26.8354
R13965 amp_biases_0.ibias3 amp_biases_0.ibias3.n7 18.7192
R13966 amp_biases_0.ibias3.n4 amp_biases_0.ibias3.t1 5.4926
R13967 amp_biases_0.ibias3.n0 amp_biases_0.ibias3.n2 4.11682
R13968 amp_biases_0.ibias3.n2 amp_biases_0.ibias3.n1 4.11576
R13969 amp_biases_0.ibias3.n3 amp_biases_0.ibias3.n1 3.20309
R13970 amp_biases_0.ibias3.n0 amp_biases_0.ibias3.n3 3.20309
R13971 amp_biases_0.ibias3.n4 amp_biases_0.ibias3.n0 2.71404
R13972 amp_biases_0.ibias3.n7 amp_biases_0.ibias3.t2 1.84683
R13973 amp_biases_0.ibias3.n7 amp_biases_0.ibias3.t3 1.84683
R13974 amp_biases_0.ibias3.n5 amp_biases_0.ibias3.n4 1.50744
R13975 amp_biases_0.ibias3.n5 amp_biases_0.ibias3.n1 1.19321
R13976 amp_biases_0.ibias3.n0 amp_biases_0.ibias3 0.953625
R13977 amp_biases_0.ibias3.n6 amp_biases_0.ibias3.n5 0.531297
R13978 amp_biases_0.ibias4.n6 amp_biases_0.ibias4.t5 281.421
R13979 amp_biases_0.ibias4.n2 amp_biases_0.ibias4.t4 232.155
R13980 amp_biases_0.ibias4.n3 amp_biases_0.ibias4.t0 232.155
R13981 amp_biases_0.ibias4 amp_biases_0.ibias4.n6 20.0327
R13982 amp_biases_0.ibias4 amp_biases_0.ibias4.n7 16.5091
R13983 amp_biases_0.ibias4.n4 amp_biases_0.ibias4.t1 5.4926
R13984 amp_biases_0.ibias4.n0 amp_biases_0.ibias4.n2 4.11682
R13985 amp_biases_0.ibias4.n2 amp_biases_0.ibias4.n1 4.11576
R13986 amp_biases_0.ibias4.n3 amp_biases_0.ibias4.n1 3.20309
R13987 amp_biases_0.ibias4.n0 amp_biases_0.ibias4.n3 3.20309
R13988 amp_biases_0.ibias4.n4 amp_biases_0.ibias4.n0 2.71404
R13989 amp_biases_0.ibias4.n7 amp_biases_0.ibias4.t2 1.84683
R13990 amp_biases_0.ibias4.n7 amp_biases_0.ibias4.t3 1.84683
R13991 amp_biases_0.ibias4.n5 amp_biases_0.ibias4.n4 1.50744
R13992 amp_biases_0.ibias4.n5 amp_biases_0.ibias4.n1 1.19321
R13993 amp_biases_0.ibias4.n0 amp_biases_0.ibias4 0.953625
R13994 amp_biases_0.ibias4.n6 amp_biases_0.ibias4.n5 0.531297
R13995 a_13231_764.n0 a_13231_764.t0 6.15493
R13996 a_13231_764.n0 a_13231_764.t2 5.15685
R13997 a_13231_764.t1 a_13231_764.n0 5.15662
R13998 a_16415_764.n0 a_16415_764.t0 6.15493
R13999 a_16415_764.n0 a_16415_764.t2 5.15685
R14000 a_16415_764.t1 a_16415_764.n0 5.15662
R14001 D83v3.n5 D83v3.n4 873.303
R14002 D83v3 D83v3.n5 585
R14003 D83v3.t1 D83v3 506.99
R14004 D83v3 D83v3.t0 150.315
R14005 D83v3.n5 D83v3.t1 147.756
R14006 D83v3.n0 D83v3.t11 104.861
R14007 D83v3.n1 D83v3.t10 104.861
R14008 D83v3.n0 D83v3.t17 104.469
R14009 D83v3.n0 D83v3.t15 104.469
R14010 D83v3.n0 D83v3.t3 104.469
R14011 D83v3.n0 D83v3.t7 104.469
R14012 D83v3.n0 D83v3.t5 104.469
R14013 D83v3.n0 D83v3.t13 104.469
R14014 D83v3.n1 D83v3.t8 104.469
R14015 D83v3.n1 D83v3.t16 104.469
R14016 D83v3.n1 D83v3.t14 104.469
R14017 D83v3.n1 D83v3.t2 104.469
R14018 D83v3.n1 D83v3.t6 104.469
R14019 D83v3.n1 D83v3.t4 104.469
R14020 D83v3.n1 D83v3.t12 104.469
R14021 D83v3.n2 D83v3.t9 99.6937
R14022 D83v3 D83v3.n3 26.513
R14023 D83v3.n0 D83v3 10.7114
R14024 D83v3.n1 D83v3 10.6036
R14025 D83v3.n2 D83v3.n0 7.19082
R14026 D83v3.n3 D83v3.n2 6.76102
R14027 D83v3.n4 D83v3 4.99562
R14028 D83v3.n3 D83v3.n1 4.65579
R14029 D83v3 D83v3.n4 2.70619
R14030 D6.n3 D6.t2 186.374
R14031 D6.n2 D6.n1 184.464
R14032 D6.n3 D6.t1 170.308
R14033 D6.n4 D6.n3 165.827
R14034 D6.n0 D6.t0 46.372
R14035 D6.n4 D6.n2 13.2781
R14036 D6.n2 D6 5.71063
R14037 D6.n1 D6 4.3525
R14038 D6 D6.n0 3.61505
R14039 D6.n0 D6 2.5677
R14040 D6.n1 D6 1.96317
R14041 D6 D6.n4 1.24229
R14042 D8.n3 D8.t1 186.374
R14043 D8.n2 D8.n1 184.464
R14044 D8.n3 D8.t0 170.308
R14045 D8.n4 D8.n3 165.827
R14046 D8.n0 D8.t2 46.372
R14047 D8.n4 D8.n2 13.2781
R14048 D8.n2 D8 5.71063
R14049 D8.n1 D8 4.3525
R14050 D8 D8.n0 3.61505
R14051 D8.n0 D8 2.5677
R14052 D8.n1 D8 1.96317
R14053 D8 D8.n4 1.24229
R14054 V1.n0 V1.t0 492.844
R14055 V1.n0 V1 13.9442
R14056 V1 V1.n0 0.063
C0 a_n2121_10269# VDD 0.902576f
C1 D83v3 a_10431_n3536# 0.042342f
C2 a_n2121_10269# a_n2603_9854# 0.024564f
C3 a_862_n8604# VDD 0.172474f
C4 a_n2559_n9065# a_n2603_n10114# 0.138963f
C5 ia_opamp_0.V2 VSS 19.0577f
C6 D13v3 a_1412_n4916# 1.31013f
C7 D03v3 AVOUT2 0.528881f
C8 D43v3 a_n1825_n338# 0.018166f
C9 a_n2577_4809# VDD 0.629385f
C10 a_n2603_7358# a_n2577_7305# 0.460789f
C11 a_n2121_7773# a_n1825_7150# 0.28899f
C12 VDD D6 0.497941f
C13 D03v3 x5.V2 0.729857f
C14 a_n2559_n9065# DVDD 0.377279f
C15 x6.V1 amp_biases_0.ibias5 0.479752f
C16 x3.R1 amp_biases_0.ibias4 0.489542f
C17 x8.V2 AVOUT2 0.613946f
C18 D53v3 VDD 1.65389f
C19 a_n2603_4862# G 0.040799f
C20 amp_biases_0.ibias1 x5.V2 0.399167f
C21 a_n2121_12765# VDD 0.870458f
C22 amp_biases_0.ibias3 amp_biases_0.ibias4 1.0136f
C23 D73v3 a_10431_n3536# 0.046327f
C24 DVDD D9 0.191057f
C25 x8.V2 x5.V2 3.06624f
C26 x3.R1 x4.V2 0.542613f
C27 a_n1825_2158# D43v3 0.17212f
C28 a_n2577_7305# VDD 0.636251f
C29 amp_biases_0.ibias3 x4.V2 1.72077f
C30 D13v3 a_n2559_8407# 0.022625f
C31 D93v3 a_10959_n3536# 0.051611f
C32 ia_opamp_0.V2 AVOUT2 1.9997f
C33 a_n2559_n6569# DVDD 0.377289f
C34 D4 V2 0.077405f
C35 D43v3 VDD 4.94409f
C36 x5.V2 ia_opamp_0.V2 0.368189f
C37 D63v3 a_10431_n3536# 0.06897f
C38 x6.V1 VOUT 2.11159f
C39 a_n2121_12765# a_n2603_12350# 0.024564f
C40 a_334_n3536# a_862_n3536# 0.104425f
C41 a_334_n3536# VSS 1.28336f
C42 a_n2559_n6569# a_n2603_n7618# 0.138963f
C43 a_10431_n8604# VSS 1.28166f
C44 D33v3 a_n1825_2158# 0.013028f
C45 a_10431_n8604# a_10959_n8604# 0.104425f
C46 a_n2577_9801# VDD 0.621838f
C47 a_n2121_10269# a_n1825_9646# 0.28899f
C48 a_1412_n9984# VDD 0.213186f
C49 D83v3 a_10959_n3536# 0.044636f
C50 a_n2603_9854# a_n2577_9801# 0.460789f
C51 a_n2559_15895# DVDD 0.377341f
C52 a_2564_12836# VSS 1.37546f
C53 a_n2121_n9699# a_n2577_n10167# 0.264713f
C54 ia_opamp_0.V2 a_1412_n4916# 0.012605f
C55 a_n2559_n4073# DVDD 0.377289f
C56 D33v3 VDD 3.24163f
C57 VDD G 0.953067f
C58 D53v3 a_10431_n3536# 0.128713f
C59 a_n2603_n10114# DVDD 0.168977f
C60 VDD D7 0.497941f
C61 ia_opamp_0.ibias VDD 5.09328f
C62 a_n1825_4654# D33v3 0.17212f
C63 a_n1825_4654# G 0.032335f
C64 a_n2577_12297# VDD 0.617081f
C65 D03v3 a_n2559_10903# 0.057171f
C66 D73v3 a_10959_n3536# 0.048324f
C67 amp_biases_0.ibias4 VDD 4.18336f
C68 x3.R1 x8.V2 0.500227f
C69 a_n2559_n1577# DVDD 0.377289f
C70 x9.V2 amp_biases_0.ibias4 4.12945f
C71 D23v3 VDD 3.11585f
C72 D93v3 a_11509_n4916# 0.458259f
C73 V2 V1 2.68736f
C74 x8.V2 amp_biases_0.ibias3 3.63465f
C75 a_n2559_15895# a_n2603_14846# 0.138963f
C76 x4.V2 VDD 9.0633f
C77 DVDD VSS 0.174825f
C78 a_n2603_n7618# DVDD 0.168977f
C79 a_n2559_n4073# a_n2603_n5122# 0.138963f
C80 VSS ibias 5.554451f
C81 x9.V2 x4.V2 0.799645f
C82 x3.R1 ia_opamp_0.V2 0.228422f
C83 a_n2121_12765# a_n1825_12142# 0.28899f
C84 a_n2603_12350# a_n2577_12297# 0.460789f
C85 D63v3 a_10959_n3536# 0.114357f
C86 a_862_n3536# VSS 1.32781f
C87 a_n2121_n7203# a_n2577_n7671# 0.264713f
C88 a_n2559_919# DVDD 0.377289f
C89 a_10959_n8604# VSS 1.32563f
C90 D13v3 VDD 3.56847f
C91 D83v3 a_11509_n4916# 0.120423f
C92 a_n2603_14846# DVDD 0.168977f
C93 a_n2121_n9699# D93v3 0.047431f
C94 a_n2603_n5122# DVDD 0.168977f
C95 a_n2559_919# VSS 0.014907f
C96 a_n1825_7150# D23v3 0.17212f
C97 AVOUT1 V2 0.012422f
C98 D53v3 a_10959_n3536# 0.592063f
C99 a_n2559_3415# DVDD 0.377289f
C100 VDD D8 0.497941f
C101 D03v3 VDD 10.3799f
C102 D73v3 a_11509_n4916# 0.163075f
C103 VSS AVOUT2 20.3182f
C104 a_n2603_n2626# DVDD 0.168977f
C105 a_n2559_3415# VSS 0.08447f
C106 a_n2559_n1577# a_n2603_n2626# 0.138963f
C107 amp_biases_0.ibias1 VDD 4.93045f
C108 x5.V2 VSS 27.2943f
C109 a_n2121_15261# a_n2577_14793# 0.264713f
C110 x8.V2 VDD 3.77323f
C111 D93v3 x6.V1 9.10921f
C112 a_n2121_n4707# a_n2577_n5175# 0.264713f
C113 a_n2559_5911# DVDD 0.377289f
C114 x9.V2 x8.V2 0.77107f
C115 D63v3 a_11509_n4916# 1.31523f
C116 a_862_n3536# a_1412_n4916# 0.19014f
C117 a_1412_n4916# VSS 1.92875f
C118 a_n2121_n7203# D83v3 0.044567f
C119 a_n2603_n130# DVDD 0.168977f
C120 a_11509_n9984# VSS 1.92492f
C121 a_10959_n8604# a_11509_n9984# 0.19014f
C122 ia_opamp_0.V2 VDD 3.02994f
C123 a_n1825_9646# D13v3 0.17212f
C124 AVOUT1 VOUT 0.100156f
C125 D83v3 x6.V1 4.89779f
C126 a_n2559_8407# DVDD 0.377289f
C127 x5.V2 AVOUT2 0.818649f
C128 a_n2559_15895# ena 0.276737f
C129 D73v3 a_n2121_n7203# 0.042392f
C130 a_n2603_2366# DVDD 0.168977f
C131 a_n2559_n9065# VDD 0.181816f
C132 a_n2559_919# a_n2603_n130# 0.138963f
C133 D03v3 a_n1825_9646# 0.010281f
C134 a_1412_n4916# AVOUT2 0.016547f
C135 x3.R1 ibias 0.022578f
C136 D73v3 x6.V1 2.58794f
C137 a_n2603_2366# VSS 0.096784f
C138 VDD D9 0.497941f
C139 a_n2121_n2211# a_n2577_n2679# 0.264713f
C140 a_n2559_10903# DVDD 0.377289f
C141 amp_biases_0.ibias2 AVOUT1 0.121094f
C142 x3.R1 VSS 23.812f
C143 a_n2121_15261# sky130_fd_sc_hvl__lsbuflv2hv_1_0[10].X 0.048684f
C144 DVDD ena 0.191399f
C145 amp_biases_0.ibias3 VSS 13.8791f
C146 a_n2121_n4707# D73v3 0.032209f
C147 a_334_n3536# VDD 0.803371f
C148 a_n2559_n6569# VDD 0.18154f
C149 D03v3 D1 0.175711f
C150 a_n2603_4862# DVDD 0.168977f
C151 a_10431_n8604# VDD 0.668038f
C152 a_n1825_12142# D03v3 0.171105f
C153 ia_opamp_0.V2 a_10431_n3536# 0.01171f
C154 D33v3 V2 0.136361f
C155 D63v3 x6.V1 1.39348f
C156 G V2 0.074334f
C157 a_n2559_13399# DVDD 0.377289f
C158 ia_opamp_0.ibias V2 0.306609f
C159 D63v3 a_n2121_n4707# 0.104034f
C160 a_n2559_15895# VDD 0.179257f
C161 a_n2603_7358# DVDD 0.168977f
C162 a_n2559_n4073# VDD 0.18218f
C163 a_n2559_3415# a_n2603_2366# 0.138963f
C164 amp_biases_0.ibias3 AVOUT2 0.112896f
C165 x3.R1 x5.V2 0.500058f
C166 D53v3 x6.V1 0.730311f
C167 D23v3 V2 0.062964f
C168 a_n2603_n10114# VDD 0.140945f
C169 a_n2121_285# a_n2577_n183# 0.264713f
C170 x4.V2 V2 0.535378f
C171 D93v3 a_334_n8604# 0.015713f
C172 amp_biases_0.ibias3 x5.V2 0.162088f
C173 amp_biases_0.ibias4 amp_biases_0.ibias5 4.71776f
C174 D13v3 D2 0.13231f
C175 D83v3 D93v3 14.5372f
C176 a_n1825_2158# VSS 0.044732f
C177 a_n2121_n2211# D63v3 0.033502f
C178 D53v3 a_n2121_n4707# 0.015263f
C179 VDD DVDD 20.706902f
C180 a_n2559_n1577# VDD 0.18154f
C181 a_n2603_9854# DVDD 0.168977f
C182 amp_biases_0.ibias5 x4.V2 2.89611f
C183 VDD ibias 0.337598f
C184 a_n2121_5277# V1 0.011508f
C185 D13v3 V2 0.062964f
C186 a_862_n3536# VDD 0.180166f
C187 x9.V2 ibias 0.017042f
C188 a_n2603_n7618# VDD 0.142356f
C189 VDD VSS 1.68051p
C190 DVDD D0 0.191057f
C191 x9.V2 VSS 21.3439f
C192 D73v3 D93v3 0.745468f
C193 D53v3 a_n2121_n2211# 0.069285f
C194 amp_biases_0.ibias4 VOUT 0.028416f
C195 a_n2603_12350# DVDD 0.168977f
C196 a_n2559_919# VDD 0.180968f
C197 a_n2559_5911# a_n2603_4862# 0.138963f
C198 AVOUT1 V1 0.406315f
C199 D03v3 V2 0.081662f
C200 D23v3 D3 0.132414f
C201 a_n2603_14846# VDD 0.142356f
C202 a_n2603_n5122# VDD 0.142356f
C203 a_n2121_2781# a_n2577_2313# 0.264713f
C204 D73v3 D83v3 10.3019f
C205 D63v3 D93v3 0.435537f
C206 VDD AVOUT2 3.43592f
C207 a_n1825_n10322# VDD 0.422564f
C208 a_n2121_285# D53v3 0.035135f
C209 D93v3 a_862_n8604# 0.012691f
C210 a_n2559_3415# VDD 0.180968f
C211 x9.V2 AVOUT2 0.381186f
C212 x5.V2 VDD 6.97056f
C213 amp_biases_0.ibias2 amp_biases_0.ibias4 0.127699f
C214 a_n2603_n2626# VDD 0.142356f
C215 x9.V2 x5.V2 0.764986f
C216 x6.V1 x4.V2 0.369149f
C217 x8.V2 amp_biases_0.ibias5 0.208521f
C218 a_10431_n3536# VSS 1.28913f
C219 a_334_n8604# a_862_n8604# 0.07931f
C220 ia_opamp_0.V2 V2 1.19672f
C221 a_n2577_4809# V1 0.011739f
C222 amp_biases_0.ibias2 x4.V2 0.228345f
C223 D53v3 D93v3 0.321343f
C224 D63v3 D83v3 0.401149f
C225 a_1412_n4916# VDD 0.20682f
C226 a_n1825_n7826# VDD 0.43082f
C227 D43v3 a_n2121_285# 0.046718f
C228 a_11509_n9984# VDD 0.016715f
C229 a_n2559_5911# VDD 0.327935f
C230 a_n2559_8407# a_n2603_7358# 0.138963f
C231 D33v3 D4 0.139956f
C232 ia_opamp_0.V2 a_11509_n4916# 0.016547f
C233 DVDD D1 0.191057f
C234 a_n2603_n130# VDD 0.142356f
C235 a_n2121_5277# a_n2577_4809# 0.264713f
C236 D63v3 D73v3 8.94018f
C237 D43v3 D93v3 0.155714f
C238 D53v3 D83v3 0.257195f
C239 a_n1825_14638# VDD 0.430705f
C240 a_n1825_n5330# VDD 0.43082f
C241 x8.V2 VOUT 0.038287f
C242 a_n2121_2781# D43v3 0.035135f
C243 a_n2559_8407# VDD 0.224805f
C244 D93v3 a_1412_n9984# 0.022752f
C245 a_n2603_2366# VDD 0.142356f
C246 D43v3 a_334_n8604# 0.049235f
C247 x3.R1 VDD 6.00188f
C248 D43v3 D5 0.146726f
C249 D43v3 D83v3 0.115078f
C250 D53v3 D73v3 0.258592f
C251 D33v3 D93v3 0.133651f
C252 a_n1825_n2834# VDD 0.43082f
C253 amp_biases_0.ibias3 VDD 5.02319f
C254 x9.V2 x3.R1 4.96863f
C255 D33v3 a_n2121_2781# 0.03444f
C256 x6.V1 x8.V2 0.367712f
C257 amp_biases_0.ibias1 amp_biases_0.ibias2 1.41657f
C258 a_n2559_10903# VDD 0.2145f
C259 a_n2559_10903# a_n2603_9854# 0.138963f
C260 a_10959_n3536# VSS 1.3278f
C261 a_n2559_n9065# a_n2121_n9699# 0.40546f
C262 x9.V2 amp_biases_0.ibias3 0.090795f
C263 D33v3 V1 0.258504f
C264 x8.V2 amp_biases_0.ibias2 0.093185f
C265 G V1 0.687566f
C266 VDD ena 0.504173f
C267 a_n2603_4862# VDD 0.191204f
C268 a_n2121_7773# a_n2577_7305# 0.264713f
C269 D33v3 a_334_n8604# 0.042342f
C270 ia_opamp_0.ibias V1 0.17087f
C271 x6.V1 ia_opamp_0.V2 0.080482f
C272 D43v3 D73v3 0.115078f
C273 D53v3 D63v3 8.48563f
C274 D33v3 D83v3 0.107562f
C275 D23v3 D93v3 0.137396f
C276 a_n1825_n338# VDD 0.43082f
C277 DVDD D2 0.191057f
C278 a_n2121_5277# D33v3 0.035135f
C279 a_n2121_5277# G 0.05594f
C280 a_n2559_13399# VDD 0.182362f
C281 D23v3 V1 0.057661f
C282 x4.V2 V1 0.324907f
C283 D53v3 D6 0.158194f
C284 a_n2603_7358# VDD 0.169958f
C285 D23v3 a_334_n8604# 0.046327f
C286 DVDD V2 0.038772f
C287 a_n2559_13399# D0 0.276737f
C288 x3.R1 a_10431_n3536# 0.31767f
C289 D43v3 D63v3 0.115078f
C290 D23v3 D83v3 0.112477f
C291 D13v3 D93v3 0.13527f
C292 D33v3 D73v3 0.107562f
C293 a_n1825_2158# VDD 0.430705f
C294 D23v3 a_n2121_5277# 0.026222f
C295 D43v3 a_862_n8604# 0.051611f
C296 a_n2559_13399# a_n2603_12350# 0.138963f
C297 VSS V2 1.61238f
C298 a_n2559_n6569# a_n2121_n7203# 0.40546f
C299 D13v3 V1 0.054525f
C300 a_n2603_9854# VDD 0.150639f
C301 a_n2121_10269# a_n2577_9801# 0.264713f
C302 a_11509_n4916# VSS 1.92882f
C303 D13v3 a_334_n8604# 0.06897f
C304 a_862_n8604# a_1412_n9984# 0.177218f
C305 a_n2121_n9699# a_n2603_n10114# 0.024564f
C306 amp_biases_0.ibias5 VSS 14.899599f
C307 x6.V1 a_10431_n8604# 0.31767f
C308 x9.V2 VDD 3.92247f
C309 D03v3 D93v3 0.199351f
C310 D23v3 D73v3 0.112477f
C311 D43v3 D53v3 1.81817f
C312 D33v3 D63v3 0.107562f
C313 D13v3 D83v3 0.111286f
C314 x4.V2 AVOUT1 1.36852f
C315 a_n1825_4654# VDD 0.431133f
C316 a_n2121_7773# D23v3 0.035135f
C317 D33v3 a_862_n8604# 0.044636f
C318 VDD D0 0.497941f
C319 a_n2121_n9699# DVDD 0.085745f
C320 D63v3 D7 0.168423f
C321 D03v3 V1 0.070054f
C322 a_n2559_10903# D1 0.276737f
C323 a_n2577_4809# G 0.045603f
C324 a_n2603_12350# VDD 0.142356f
C325 D03v3 a_334_n8604# 0.164977f
C326 amp_biases_0.ibias1 V1 0.320387f
C327 DVDD D3 0.191057f
C328 a_n2559_3415# V2 0.01892f
C329 D13v3 D73v3 0.111286f
C330 D33v3 D53v3 0.123472f
C331 D23v3 D63v3 0.112477f
C332 D03v3 D83v3 0.118929f
C333 a_n1825_7150# VDD 0.468134f
C334 D13v3 a_n2121_7773# 0.021443f
C335 D23v3 a_862_n8604# 0.048325f
C336 VSS VOUT 16.3614f
C337 a_n2559_15895# a_n2121_15261# 0.40546f
C338 a_n2121_n7203# DVDD 0.085745f
C339 D93v3 ia_opamp_0.V2 0.970198f
C340 a_n2559_n4073# a_n2121_n4707# 0.40546f
C341 x3.R1 a_10959_n3536# 0.145098f
C342 amp_biases_0.ibias5 x5.V2 0.118815f
C343 D43v3 a_1412_n9984# 0.458259f
C344 a_n2121_12765# a_n2577_12297# 0.264713f
C345 a_10431_n3536# VDD 0.651327f
C346 ia_opamp_0.V2 V1 0.302013f
C347 a_n2121_n7203# a_n2603_n7618# 0.024564f
C348 D03v3 AVOUT1 0.024603f
C349 x6.V1 ibias 0.016798f
C350 D73v3 D8 0.167459f
C351 D03v3 D73v3 0.117069f
C352 D23v3 D53v3 0.128352f
C353 D13v3 D63v3 0.111286f
C354 D33v3 D43v3 11.4682f
C355 a_n1825_9646# VDD 0.447291f
C356 a_n2121_10269# D13v3 0.034184f
C357 D13v3 a_862_n8604# 0.140391f
C358 a_n2559_8407# D2 0.276737f
C359 amp_biases_0.ibias1 AVOUT1 3.22644f
C360 a_n2603_n10114# a_n2577_n10167# 0.460789f
C361 a_n2559_n9065# D93v3 0.015265f
C362 x6.V1 VSS 32.8241f
C363 a_n2121_n9699# a_n1825_n10322# 0.28899f
C364 a_n2121_15261# DVDD 0.085745f
C365 x6.V1 a_10959_n8604# 0.154322f
C366 a_n2121_n4707# DVDD 0.085745f
C367 D83v3 ia_opamp_0.V2 0.789011f
C368 x8.V2 AVOUT1 0.377184f
C369 amp_biases_0.ibias2 VSS 13.3701f
C370 D33v3 a_1412_n9984# 0.120423f
C371 AVOUT2 VOUT 0.174328f
C372 a_n2577_n10167# DVDD 0.103609f
C373 VDD D1 0.516651f
C374 D23v3 D43v3 0.616188f
C375 D13v3 D53v3 0.127141f
C376 D03v3 D63v3 0.117035f
C377 D33v3 G 0.018841f
C378 a_n1825_12142# VDD 0.431406f
C379 D43v3 x4.V2 9.14715f
C380 D03v3 a_n2121_10269# 0.094739f
C381 D03v3 a_862_n8604# 1.046f
C382 ia_opamp_0.V2 AVOUT1 0.986075f
C383 D73v3 ia_opamp_0.V2 0.670971f
C384 D93v3 a_10431_n8604# 0.061799f
C385 a_n2121_n2211# DVDD 0.085745f
C386 a_n2559_n1577# a_n2121_n2211# 0.40546f
C387 DVDD D4 0.191057f
C388 D23v3 a_1412_n9984# 0.20376f
C389 a_n2121_15261# a_n2603_14846# 0.024564f
C390 D83v3 D9 0.122407f
C391 a_n2577_n7671# DVDD 0.103827f
C392 a_n2121_n4707# a_n2603_n5122# 0.024564f
C393 x3.R1 a_11509_n4916# 0.710767f
C394 a_n2559_5911# D3 0.276737f
C395 amp_biases_0.ibias2 AVOUT2 3.25165f
C396 VSS D4 0.036767f
C397 D13v3 D43v3 0.307857f
C398 x6.V1 x5.V2 0.372989f
C399 D03v3 D53v3 0.132881f
C400 D23v3 D33v3 9.03536f
C401 x3.R1 amp_biases_0.ibias5 0.130422f
C402 D23v3 G 0.086867f
C403 a_n2121_12765# D03v3 0.03394f
C404 D33v3 x4.V2 5.01902f
C405 a_n2603_n7618# a_n2577_n7671# 0.460789f
C406 a_n2121_n7203# a_n1825_n7826# 0.28899f
C407 amp_biases_0.ibias2 x5.V2 0.248886f
C408 amp_biases_0.ibias3 amp_biases_0.ibias5 0.135327f
C409 D83v3 a_10431_n8604# 0.042342f
C410 a_n2121_285# DVDD 0.085745f
C411 D63v3 ia_opamp_0.V2 0.610716f
C412 ia_opamp_0.ibias x4.V2 0.130926f
C413 D13v3 a_1412_n9984# 1.72752f
C414 a_n2577_14793# DVDD 0.103827f
C415 a_n2577_n5175# DVDD 0.103827f
C416 amp_biases_0.ibias4 x4.V2 2.33031f
C417 x6.V1 a_11509_n9984# 0.710767f
C418 D03v3 D43v3 0.192773f
C419 D13v3 D33v3 0.289863f
C420 D13v3 G 0.066858f
C421 D23v3 x4.V2 2.71456f
C422 D73v3 a_n2559_n6569# 0.04344f
C423 D53v3 ia_opamp_0.V2 0.656723f
C424 a_n2121_2781# DVDD 0.085745f
C425 D73v3 a_10431_n8604# 0.046327f
C426 x3.R1 VOUT 0.58027f
C427 a_n2559_919# a_n2121_285# 0.40546f
C428 a_n2559_3415# D4 0.276737f
C429 VDD D2 0.515529f
C430 DVDD V1 0.029725f
C431 sky130_fd_sc_hvl__lsbuflv2hv_1_0[10].X a_2564_12836# 1.41702f
C432 amp_biases_0.ibias3 VOUT 0.026535f
C433 D93v3 VSS 21.358f
C434 D93v3 a_10959_n8604# 0.064191f
C435 a_n2577_n2679# DVDD 0.103827f
C436 a_n2121_2781# VSS 0.187137f
C437 a_n2121_n2211# a_n2603_n2626# 0.024564f
C438 D03v3 D33v3 0.145037f
C439 D13v3 D23v3 8.33479f
C440 D03v3 G 0.139181f
C441 a_n2121_15261# a_n1825_14638# 0.28899f
C442 VSS V1 1.1636f
C443 a_n2603_14846# a_n2577_14793# 0.460789f
C444 a_n2559_15895# sky130_fd_sc_hvl__lsbuflv2hv_1_0[10].X 0.01643f
C445 D13v3 x4.V2 1.52523f
C446 DVDD D5 0.191057f
C447 VDD V2 0.596698f
C448 a_n2603_n5122# a_n2577_n5175# 0.460789f
C449 a_n2121_n4707# a_n1825_n5330# 0.28899f
C450 D43v3 ia_opamp_0.V2 0.487025f
C451 D63v3 a_10431_n8604# 0.069056f
C452 a_n2121_5277# DVDD 0.085745f
C453 a_10431_n3536# a_10959_n3536# 0.104425f
C454 D03v3 ia_opamp_0.ibias 0.080425f
C455 a_334_n8604# VSS 1.27872f
C456 x6.V1 x3.R1 0.655356f
C457 VSS D5 0.017931f
C458 D83v3 VSS 13.590401f
C459 D83v3 a_10959_n8604# 0.044636f
C460 a_n2577_n183# DVDD 0.103827f
C461 ia_opamp_0.ibias amp_biases_0.ibias1 0.888026f
C462 amp_biases_0.ibias5 VDD 4.13942f
C463 D03v3 D23v3 0.146354f
C464 amp_biases_0.ibias1 amp_biases_0.ibias4 0.035418f
C465 amp_biases_0.ibias2 amp_biases_0.ibias3 2.55697f
C466 D03v3 x4.V2 0.958425f
C467 x9.V2 amp_biases_0.ibias5 0.345488f
C468 a_n1825_n10322# D93v3 0.177675f
C469 a_n2559_919# D5 0.276737f
C470 x8.V2 amp_biases_0.ibias4 0.256731f
C471 D63v3 a_n2559_n4073# 0.049556f
C472 sky130_fd_sc_hvl__lsbuflv2hv_1_0[10].X ibias 1.86202f
C473 a_n2121_7773# DVDD 0.085745f
C474 D53v3 a_10431_n8604# 0.163876f
C475 D33v3 ia_opamp_0.V2 0.421775f
C476 a_n2559_3415# a_n2121_2781# 0.40546f
C477 ia_opamp_0.V2 G 0.284326f
C478 D93v3 x5.V2 0.129642f
C479 amp_biases_0.ibias1 x4.V2 0.274329f
C480 VSS AVOUT1 18.336f
C481 sky130_fd_sc_hvl__lsbuflv2hv_1_0[10].X VSS 4.56822f
C482 x8.V2 x4.V2 0.781675f
C483 D73v3 VSS 9.8428f
C484 ia_opamp_0.ibias ia_opamp_0.V2 4.0119f
C485 a_n2577_2313# DVDD 0.103827f
C486 a_n2121_n9699# VDD 0.866649f
C487 D73v3 a_10959_n8604# 0.048347f
C488 a_n2121_285# a_n2603_n130# 0.024564f
C489 x5.V2 V1 0.359942f
C490 D03v3 D13v3 8.298651f
C491 x5.V2 a_334_n8604# 0.31767f
C492 D43v3 a_334_n3536# 0.049251f
C493 VDD VOUT 2.93085f
C494 D93v3 a_11509_n9984# 0.481011f
C495 a_n2577_2313# VSS 0.091931f
C496 a_n2603_n2626# a_n2577_n2679# 0.460789f
C497 a_n2121_n2211# a_n1825_n2834# 0.28899f
C498 VDD D3 0.970763f
C499 a_n2121_10269# DVDD 0.085745f
C500 D23v3 ia_opamp_0.V2 0.343735f
C501 D83v3 x5.V2 0.103819f
C502 x4.V2 ia_opamp_0.V2 2.44294f
C503 x9.V2 VOUT 0.061359f
C504 D63v3 VSS 7.24861f
C505 D63v3 a_10959_n8604# 0.130644f
C506 a_n2577_4809# DVDD 0.103827f
C507 a_n2121_n7203# VDD 0.86946f
C508 DVDD D6 0.191057f
C509 a_862_n8604# VSS 1.27579f
C510 a_n2559_n1577# D6 0.276737f
C511 AVOUT1 AVOUT2 1.58936f
C512 a_n1825_n7826# D83v3 0.179047f
C513 x6.V1 VDD 7.84011f
C514 D83v3 a_11509_n9984# 0.120423f
C515 D33v3 a_334_n3536# 0.042361f
C516 D53v3 a_n2559_n1577# 0.043381f
C517 a_n2121_12765# DVDD 0.085745f
C518 x5.V2 AVOUT1 3.22467f
C519 D13v3 ia_opamp_0.V2 0.012164f
C520 a_n2559_5911# a_n2121_5277# 0.40546f
C521 D73v3 x5.V2 0.103819f
C522 x6.V1 x9.V2 0.471563f
C523 amp_biases_0.ibias2 VDD 5.04202f
C524 D53v3 VSS 7.23672f
C525 a_n2121_15261# VDD 0.869226f
C526 a_n2577_7305# DVDD 0.103827f
C527 a_n2121_n4707# VDD 0.86946f
C528 D53v3 a_10959_n8604# 0.979915f
C529 a_n2121_2781# a_n2603_2366# 0.024564f
C530 D93v3 x3.R1 9.16655f
C531 D23v3 a_334_n3536# 0.046349f
C532 a_n2577_n10167# VDD 0.602952f
C533 D73v3 a_11509_n9984# 0.18595f
C534 a_n2603_n130# a_n2577_n183# 0.460789f
C535 a_n2121_285# a_n1825_n338# 0.28899f
C536 x4.V2 a_334_n3536# 0.369513f
C537 D03v3 ia_opamp_0.V2 0.067993f
C538 D63v3 x5.V2 0.103819f
C539 x5.V2 a_862_n8604# 0.154322f
C540 a_n2559_n4073# D7 0.276737f
C541 D43v3 a_862_n3536# 0.051611f
C542 D43v3 VSS 13.219901f
C543 a_n2121_n2211# VDD 0.86946f
C544 a_n2577_9801# DVDD 0.103827f
C545 D83v3 x3.R1 4.91473f
C546 VDD D4 0.497941f
C547 a_n1825_14638# sky130_fd_sc_hvl__lsbuflv2hv_1_0[10].X 0.17815f
C548 D53v3 AVOUT2 0.579576f
C549 a_n1825_n5330# D73v3 0.16854f
C550 a_n2577_n7671# VDD 0.617081f
C551 D63v3 a_11509_n9984# 1.7019f
C552 D13v3 a_334_n3536# 0.069018f
C553 DVDD G 0.04073f
C554 D43v3 a_n2559_919# 0.035884f
C555 a_10959_n3536# a_11509_n4916# 0.19014f
C556 a_1412_n9984# VSS 1.89089f
C557 a_n2559_8407# a_n2121_7773# 0.40546f
C558 D53v3 x5.V2 0.118754f
C559 DVDD D7 0.191057f
C560 D33v3 a_862_n3536# 0.044636f
C561 D33v3 VSS 8.37378f
C562 VSS G 1.26683f
C563 a_n2577_12297# DVDD 0.103827f
C564 a_n2121_285# VDD 0.869345f
C565 a_n2121_5277# a_n2603_4862# 0.024564f
C566 D73v3 x3.R1 2.60579f
C567 D43v3 AVOUT2 1.12907f
C568 ia_opamp_0.ibias VSS 12.9859f
C569 D63v3 a_n1825_n5330# 0.043534f
C570 a_n2577_14793# VDD 0.617081f
C571 D03v3 a_334_n3536# 0.098881f
C572 a_n2577_n5175# VDD 0.617081f
C573 a_n2603_2366# a_n2577_2313# 0.460789f
C574 a_n2559_n6569# D8 0.276737f
C575 a_n2121_2781# a_n1825_2158# 0.28899f
C576 amp_biases_0.ibias4 VSS 13.594299f
C577 D43v3 x5.V2 9.157269f
C578 D23v3 a_862_n3536# 0.048324f
C579 D93v3 VDD 2.6743f
C580 D23v3 VSS 5.04317f
C581 x4.V2 a_862_n3536# 0.154411f
C582 a_n2121_2781# VDD 0.869226f
C583 x4.V2 VSS 27.193699f
C584 D63v3 x3.R1 1.41646f
C585 x5.V2 a_1412_n9984# 0.710781f
C586 D43v3 a_1412_n4916# 0.458259f
C587 VDD V1 2.84542f
C588 D33v3 AVOUT2 0.704691f
C589 a_n1825_n2834# D63v3 0.169603f
C590 a_n2577_n2679# VDD 0.617081f
C591 D33v3 a_n2559_3415# 0.029984f
C592 a_334_n8604# VDD 0.849494f
C593 a_n2559_10903# a_n2121_10269# 0.40546f
C594 D33v3 x5.V2 6.02239f
C595 a_n1825_4654# V1 0.024216f
C596 D13v3 a_862_n3536# 0.102325f
C597 VDD D5 0.497941f
C598 D83v3 VDD 1.10488f
C599 D13v3 VSS 3.32471f
C600 a_n2121_5277# VDD 0.958818f
C601 a_n2121_7773# a_n2603_7358# 0.024564f
C602 D53v3 x3.R1 0.793176f
C603 a_n2559_n9065# D9 0.276737f
C604 amp_biases_0.ibias4 x5.V2 0.111193f
C605 D33v3 a_1412_n4916# 0.120423f
C606 D23v3 AVOUT2 0.61129f
C607 D53v3 a_n1825_n2834# 0.027586f
C608 x4.V2 AVOUT2 0.333907f
C609 DVDD D8 0.191057f
C610 a_n2577_n183# VDD 0.617081f
C611 a_n2603_4862# a_n2577_4809# 0.460789f
C612 a_n2121_5277# a_n1825_4654# 0.28899f
C613 D23v3 x5.V2 2.7691f
C614 x5.V2 x4.V2 0.702101f
C615 sky130_fd_sc_hvl__lsbuflv2hv_1_0[10].X VDD 1.1285f
C616 VDD AVOUT1 3.19587f
C617 D03v3 a_862_n3536# 0.561931f
C618 D73v3 VDD 0.971707f
C619 D03v3 VSS 3.44989f
C620 a_n2121_7773# VDD 0.924078f
C621 D93v3 a_10431_n3536# 0.049235f
C622 x8.V2 ibias 0.012661f
C623 amp_biases_0.ibias1 VSS 12.997201f
C624 D13v3 AVOUT2 0.553347f
C625 D23v3 a_1412_n4916# 0.156861f
C626 a_n1825_n338# D53v3 0.17212f
C627 sky130_fd_sc_hvl__lsbuflv2hv_1_0[10].X D0 0.122407f
C628 x4.V2 a_1412_n4916# 0.710811f
C629 a_n2577_2313# VDD 0.617081f
C630 x8.V2 VSS 20.8212f
C631 D23v3 a_n2559_5911# 0.024032f
C632 a_n2559_13399# a_n2121_12765# 0.40546f
C633 D13v3 x5.V2 1.38312f
C634 amp_biases_0.ibias5 VOUT 2.95501f
C635 D63v3 VDD 0.978429f
C636 V1 DVSS 3.132558f
C637 V2 DVSS 1.70795f
C638 G DVSS 0.62531f
C639 VOUT DVSS 7.264884f
C640 AVOUT2 DVSS 7.541774f
C641 AVOUT1 DVSS 7.016088f
C642 ibias DVSS 5.69287f
C643 D9 DVSS 1.2133f
C644 D8 DVSS 1.21022f
C645 D7 DVSS 1.20998f
C646 D6 DVSS 1.21033f
C647 D5 DVSS 1.21045f
C648 D4 DVSS 1.21057f
C649 D3 DVSS 1.2083f
C650 D2 DVSS 1.21084f
C651 D1 DVSS 1.20986f
C652 D0 DVSS 1.2133f
C653 ena DVSS 1.31678f
C654 VSS DVSS 57.050907f
C655 DVDD DVSS 16.149006f
C656 VDD DVSS 2.122794p
C657 a_11509_n9984# DVSS 0.459944f
C658 a_10959_n8604# DVSS 0.229403f
C659 a_10431_n8604# DVSS 0.229036f
C660 a_1412_n9984# DVSS 0.463242f
C661 a_862_n8604# DVSS 0.229373f
C662 a_334_n8604# DVSS 0.229036f
C663 a_11509_n4916# DVSS 0.479204f
C664 a_10959_n3536# DVSS 0.23607f
C665 a_10431_n3536# DVSS 0.239515f
C666 a_1412_n4916# DVSS 0.482503f
C667 a_862_n3536# DVSS 0.239867f
C668 a_334_n3536# DVSS 0.239515f
C669 ia_opamp_0.V2 DVSS 8.417559f
C670 x4.V2 DVSS 10.900803f
C671 x5.V2 DVSS 9.615119f
C672 amp_biases_0.ibias5 DVSS 12.50264f
C673 amp_biases_0.ibias4 DVSS 10.826969f
C674 amp_biases_0.ibias3 DVSS 7.494782f
C675 amp_biases_0.ibias2 DVSS 6.50279f
C676 amp_biases_0.ibias1 DVSS 5.825887f
C677 ia_opamp_0.ibias DVSS 6.141258f
C678 x8.V2 DVSS 8.113983f
C679 x3.R1 DVSS 9.157716f
C680 x9.V2 DVSS 8.230323f
C681 x6.V1 DVSS 10.166674f
C682 a_2564_12836# DVSS 0.418398f
C683 D93v3 DVSS 15.803851f
C684 a_n1825_n10322# DVSS 0.508832f
C685 a_n2577_n10167# DVSS 0.891524f
C686 a_n2603_n10114# DVSS 1.7004f
C687 a_n2121_n9699# DVSS 1.53725f
C688 a_n2559_n9065# DVSS 1.95881f
C689 D83v3 DVSS 11.389816f
C690 a_n1825_n7826# DVSS 0.502625f
C691 a_n2577_n7671# DVSS 0.869809f
C692 a_n2603_n7618# DVSS 1.69935f
C693 a_n2121_n7203# DVSS 1.53217f
C694 a_n2559_n6569# DVSS 1.95873f
C695 D73v3 DVSS 9.83117f
C696 a_n1825_n5330# DVSS 0.502625f
C697 a_n2577_n5175# DVSS 0.869809f
C698 a_n2603_n5122# DVSS 1.69935f
C699 a_n2121_n4707# DVSS 1.53217f
C700 a_n2559_n4073# DVSS 1.95873f
C701 D63v3 DVSS 8.857109f
C702 a_n1825_n2834# DVSS 0.502625f
C703 a_n2577_n2679# DVSS 0.869809f
C704 a_n2603_n2626# DVSS 1.69935f
C705 a_n2121_n2211# DVSS 1.53217f
C706 a_n2559_n1577# DVSS 1.95873f
C707 D53v3 DVSS 9.894689f
C708 a_n1825_n338# DVSS 0.502625f
C709 a_n2577_n183# DVSS 0.869809f
C710 a_n2603_n130# DVSS 1.69935f
C711 a_n2121_285# DVSS 1.53217f
C712 a_n2559_919# DVSS 1.95846f
C713 D43v3 DVSS 14.41423f
C714 a_n1825_2158# DVSS 0.502625f
C715 a_n2577_2313# DVSS 0.869809f
C716 a_n2603_2366# DVSS 1.69935f
C717 a_n2121_2781# DVSS 1.53217f
C718 a_n2559_3415# DVSS 1.95873f
C719 D33v3 DVSS 12.386173f
C720 a_n1825_4654# DVSS 0.501931f
C721 a_n2577_4809# DVSS 0.869809f
C722 a_n2603_4862# DVSS 1.69935f
C723 a_n2121_5277# DVSS 1.53217f
C724 a_n2559_5911# DVSS 1.95873f
C725 D23v3 DVSS 11.655425f
C726 a_n1825_7150# DVSS 0.502625f
C727 a_n2577_7305# DVSS 0.869809f
C728 a_n2603_7358# DVSS 1.69935f
C729 a_n2121_7773# DVSS 1.53217f
C730 a_n2559_8407# DVSS 1.95873f
C731 D13v3 DVSS 10.486039f
C732 a_n1825_9646# DVSS 0.502625f
C733 a_n2577_9801# DVSS 0.869809f
C734 a_n2603_9854# DVSS 1.69935f
C735 a_n2121_10269# DVSS 1.53217f
C736 a_n2559_10903# DVSS 1.95873f
C737 D03v3 DVSS 13.179908f
C738 a_n1825_12142# DVSS 0.50249f
C739 a_n2577_12297# DVSS 0.869809f
C740 a_n2603_12350# DVSS 1.69935f
C741 a_n2121_12765# DVSS 1.53217f
C742 a_n2559_13399# DVSS 1.95873f
C743 sky130_fd_sc_hvl__lsbuflv2hv_1_0[10].X DVSS 2.548698f
C744 a_n1825_14638# DVSS 0.502625f
C745 a_n2577_14793# DVSS 0.869809f
C746 a_n2603_14846# DVSS 1.69981f
C747 a_n2121_15261# DVSS 1.53427f
C748 a_n2559_15895# DVSS 1.96945f
C749 V1.t0 DVSS 1.36383f
C750 V1.n0 DVSS 1.68341f
C751 D83v3.n0 DVSS 11.9775f
C752 D83v3.n1 DVSS 14.3103f
C753 D83v3.t0 DVSS 0.045073f
C754 D83v3.t9 DVSS 0.952299f
C755 D83v3.t11 DVSS 1.02051f
C756 D83v3.t13 DVSS 1.0151f
C757 D83v3.t5 DVSS 1.0151f
C758 D83v3.t7 DVSS 1.0151f
C759 D83v3.t3 DVSS 1.0151f
C760 D83v3.t15 DVSS 1.0151f
C761 D83v3.t17 DVSS 1.0151f
C762 D83v3.n2 DVSS 1.62591f
C763 D83v3.t10 DVSS 1.02051f
C764 D83v3.t12 DVSS 1.0151f
C765 D83v3.t4 DVSS 1.0151f
C766 D83v3.t6 DVSS 1.0151f
C767 D83v3.t2 DVSS 1.0151f
C768 D83v3.t14 DVSS 1.0151f
C769 D83v3.t16 DVSS 1.0151f
C770 D83v3.t8 DVSS 1.01506f
C771 D83v3.n3 DVSS 6.37411f
C772 D83v3.n4 DVSS 0.038015f
C773 D83v3.t1 DVSS 0.042327f
C774 D83v3.n5 DVSS 0.037338f
C775 a_16415_764.t0 DVSS 1.02739f
C776 a_16415_764.t2 DVSS 0.830152f
C777 a_16415_764.n0 DVSS 7.41434f
C778 a_16415_764.t1 DVSS 0.828116f
C779 a_13231_764.t0 DVSS 1.31221f
C780 a_13231_764.t2 DVSS 1.06029f
C781 a_13231_764.n0 DVSS 9.4698f
C782 a_13231_764.t1 DVSS 1.05769f
C783 amp_biases_0.ibias4.n0 DVSS 2.49894f
C784 amp_biases_0.ibias4.n1 DVSS 2.17573f
C785 amp_biases_0.ibias4.t4 DVSS 2.17682f
C786 amp_biases_0.ibias4.n2 DVSS 2.29498f
C787 amp_biases_0.ibias4.t0 DVSS 2.17682f
C788 amp_biases_0.ibias4.n3 DVSS 1.77993f
C789 amp_biases_0.ibias4.t1 DVSS 0.937854f
C790 amp_biases_0.ibias4.n4 DVSS 2.48805f
C791 amp_biases_0.ibias4.n5 DVSS 0.587334f
C792 amp_biases_0.ibias4.t5 DVSS 2.68616f
C793 amp_biases_0.ibias4.n6 DVSS 7.87514f
C794 amp_biases_0.ibias4.t2 DVSS 0.250794f
C795 amp_biases_0.ibias4.t3 DVSS 0.250794f
C796 amp_biases_0.ibias4.n7 DVSS 0.999407f
C797 amp_biases_0.ibias3.n0 DVSS 2.19883f
C798 amp_biases_0.ibias3.n1 DVSS 1.91444f
C799 amp_biases_0.ibias3.t4 DVSS 1.91539f
C800 amp_biases_0.ibias3.n2 DVSS 2.01937f
C801 amp_biases_0.ibias3.t0 DVSS 1.91539f
C802 amp_biases_0.ibias3.n3 DVSS 1.56617f
C803 amp_biases_0.ibias3.t1 DVSS 0.825223f
C804 amp_biases_0.ibias3.n4 DVSS 2.18925f
C805 amp_biases_0.ibias3.n5 DVSS 0.516798f
C806 amp_biases_0.ibias3.t5 DVSS 2.36357f
C807 amp_biases_0.ibias3.n6 DVSS 7.16947f
C808 amp_biases_0.ibias3.t2 DVSS 0.220675f
C809 amp_biases_0.ibias3.t3 DVSS 0.220675f
C810 amp_biases_0.ibias3.n7 DVSS 1.18911f
C811 a_9782_281.t1 DVSS 4.66674f
C812 a_9782_281.t0 DVSS 0.133257f
C813 a_12966_281.t1 DVSS 4.66674f
C814 a_12966_281.t0 DVSS 0.133257f
C815 ibias.t0 DVSS 0.961891f
C816 a_2622_12748.t0 DVSS 0.169392f
C817 a_2622_12748.t1 DVSS 1.43945f
C818 a_2622_12748.t3 DVSS 1.44644f
C819 a_2622_12748.n0 DVSS 4.40059f
C820 a_2622_12748.n1 DVSS 0.57474f
C821 a_2622_12748.t2 DVSS 0.169392f
C822 sky130_fd_sc_hvl__lsbuflv2hv_1_0[10].X.t0 DVSS 0.013087f
C823 sky130_fd_sc_hvl__lsbuflv2hv_1_0[10].X.t2 DVSS 0.73596f
C824 sky130_fd_sc_hvl__lsbuflv2hv_1_0[10].X.t3 DVSS 0.732087f
C825 sky130_fd_sc_hvl__lsbuflv2hv_1_0[10].X.n0 DVSS 2.26174f
C826 sky130_fd_sc_hvl__lsbuflv2hv_1_0[10].X.n1 DVSS 0.011038f
C827 sky130_fd_sc_hvl__lsbuflv2hv_1_0[10].X.t1 DVSS 0.01229f
C828 sky130_fd_sc_hvl__lsbuflv2hv_1_0[10].X.n2 DVSS 0.010841f
C829 a_6598_281.t1 DVSS 4.66674f
C830 a_6598_281.t0 DVSS 0.133257f
C831 a_6863_764.t0 DVSS 1.00705f
C832 a_6863_764.t2 DVSS 0.811718f
C833 a_6863_764.n0 DVSS 7.26752f
C834 a_6863_764.t1 DVSS 0.813714f
C835 a_13767_764.t0 DVSS 0.18974f
C836 a_13767_764.n0 DVSS 1.1588f
C837 a_13767_764.n1 DVSS 3.40015f
C838 a_13767_764.t7 DVSS 1.97165f
C839 a_13767_764.n2 DVSS 0.473297f
C840 a_13767_764.t6 DVSS 1.97165f
C841 a_13767_764.n3 DVSS 0.015846f
C842 a_13767_764.n4 DVSS 3.4092f
C843 a_13767_764.n5 DVSS 1.86827f
C844 a_13767_764.t4 DVSS 1.97165f
C845 a_13767_764.n6 DVSS 0.016627f
C846 a_13767_764.n7 DVSS 1.86628f
C847 a_13767_764.t5 DVSS 1.97165f
C848 a_13767_764.n8 DVSS 1.53199f
C849 a_13767_764.n9 DVSS 1.05306f
C850 a_13767_764.t2 DVSS 10.505401f
C851 a_13767_764.n10 DVSS 0.853045f
C852 a_13767_764.t3 DVSS 1.64215f
C853 a_13767_764.n11 DVSS 1.45288f
C854 a_13767_764.n12 DVSS 0.386963f
C855 a_13767_764.t1 DVSS 0.18974f
C856 a_3414_281.t1 DVSS 4.66674f
C857 a_3414_281.t0 DVSS 0.133257f
C858 amp_biases_0.ibias2.n0 DVSS 2.18148f
C859 amp_biases_0.ibias2.n1 DVSS 1.89933f
C860 amp_biases_0.ibias2.t4 DVSS 1.90028f
C861 amp_biases_0.ibias2.n2 DVSS 2.00343f
C862 amp_biases_0.ibias2.t0 DVSS 1.90028f
C863 amp_biases_0.ibias2.n3 DVSS 1.55381f
C864 amp_biases_0.ibias2.t1 DVSS 0.818712f
C865 amp_biases_0.ibias2.n4 DVSS 2.17198f
C866 amp_biases_0.ibias2.n5 DVSS 0.512721f
C867 amp_biases_0.ibias2.t5 DVSS 2.34492f
C868 amp_biases_0.ibias2.n6 DVSS 6.51229f
C869 amp_biases_0.ibias2.t3 DVSS 0.218934f
C870 amp_biases_0.ibias2.t2 DVSS 0.218934f
C871 amp_biases_0.ibias2.n7 DVSS 1.34931f
C872 a_2308_n4916.t3 DVSS 0.198045f
C873 a_2308_n4916.t2 DVSS 0.043897f
C874 a_2308_n4916.t1 DVSS 0.043897f
C875 a_2308_n4916.n0 DVSS 0.127895f
C876 a_2308_n4916.n1 DVSS 0.534999f
C877 a_2308_n4916.t0 DVSS 0.1543f
C878 a_2308_n4916.n2 DVSS 0.372322f
C879 a_2308_n4916.t6 DVSS 0.067673f
C880 a_2308_n4916.t5 DVSS 0.065867f
C881 a_2308_n4916.n3 DVSS 1.20595f
C882 a_2308_n4916.t7 DVSS 0.065867f
C883 a_2308_n4916.n4 DVSS 0.643717f
C884 a_2308_n4916.n5 DVSS 0.78373f
C885 a_2308_n4916.t4 DVSS 0.291836f
C886 a_2308_n9984.t3 DVSS 0.215267f
C887 a_2308_n9984.t2 DVSS 0.047715f
C888 a_2308_n9984.t1 DVSS 0.047715f
C889 a_2308_n9984.n0 DVSS 0.139017f
C890 a_2308_n9984.n1 DVSS 0.581521f
C891 a_2308_n9984.t0 DVSS 0.167717f
C892 a_2308_n9984.n2 DVSS 0.404698f
C893 a_2308_n9984.t6 DVSS 0.073558f
C894 a_2308_n9984.t7 DVSS 0.071595f
C895 a_2308_n9984.n3 DVSS 1.31082f
C896 a_2308_n9984.t5 DVSS 0.071595f
C897 a_2308_n9984.n4 DVSS 0.699693f
C898 a_2308_n9984.n5 DVSS 0.851881f
C899 a_2308_n9984.t4 DVSS 0.317213f
C900 D23v3.n0 DVSS 5.76463f
C901 D23v3.n1 DVSS 6.21323f
C902 D23v3.t0 DVSS 0.049363f
C903 D23v3.t9 DVSS 1.16123f
C904 D23v3.t5 DVSS 1.1553f
C905 D23v3.t7 DVSS 1.15526f
C906 D23v3.t3 DVSS 1.08666f
C907 D23v3.t2 DVSS 1.0883f
C908 D23v3.t8 DVSS 1.16123f
C909 D23v3.t4 DVSS 1.1553f
C910 D23v3.t6 DVSS 1.15526f
C911 D23v3.n2 DVSS 3.69958f
C912 D23v3.n3 DVSS 3.40527f
C913 D23v3.n4 DVSS 0.041634f
C914 D23v3.t1 DVSS 0.046357f
C915 D23v3.n5 DVSS 0.040892f
C916 amp_biases_0.ibias5.n0 DVSS 2.40913f
C917 amp_biases_0.ibias5.n1 DVSS 5.49715f
C918 amp_biases_0.ibias5.t4 DVSS 2.59853f
C919 amp_biases_0.ibias5.t5 DVSS 2.09858f
C920 amp_biases_0.ibias5.n2 DVSS 2.2125f
C921 amp_biases_0.ibias5.t0 DVSS 2.09858f
C922 amp_biases_0.ibias5.n3 DVSS 1.71596f
C923 amp_biases_0.ibias5.t1 DVSS 0.904147f
C924 amp_biases_0.ibias5.n4 DVSS 2.39912f
C925 amp_biases_0.ibias5.n5 DVSS 5.32003f
C926 amp_biases_0.ibias5.t3 DVSS 0.241781f
C927 amp_biases_0.ibias5.t2 DVSS 0.241781f
C928 amp_biases_0.ibias5.n6 DVSS 0.859542f
C929 D13v3.n0 DVSS 2.06728f
C930 D13v3.t0 DVSS 0.045901f
C931 D13v3.t3 DVSS 1.11425f
C932 D13v3.t5 DVSS 1.04338f
C933 D13v3.t4 DVSS 1.04553f
C934 D13v3.t2 DVSS 1.11425f
C935 D13v3.n1 DVSS 2.39235f
C936 D13v3.n2 DVSS 3.4941f
C937 D13v3.n3 DVSS 3.19868f
C938 D13v3.n4 DVSS 0.038714f
C939 D13v3.t1 DVSS 0.043105f
C940 D13v3.n5 DVSS 0.038024f
C941 D53v3.n0 DVSS 6.4941f
C942 D53v3.t0 DVSS 0.035289f
C943 D53v3.t3 DVSS 0.792256f
C944 D53v3.n1 DVSS 1.49389f
C945 D53v3.t2 DVSS 0.840693f
C946 D53v3.n2 DVSS 0.029763f
C947 D53v3.t1 DVSS 0.03314f
C948 D53v3.n3 DVSS 0.029233f
C949 a_3679_764.t0 DVSS 0.986702f
C950 a_3679_764.t2 DVSS 0.797275f
C951 a_3679_764.n0 DVSS 7.1207f
C952 a_3679_764.t1 DVSS 0.795319f
C953 V2.t0 DVSS 0.792874f
C954 V2.n0 DVSS 0.8022f
C955 a_7399_764.t0 DVSS 0.17422f
C956 a_7399_764.n0 DVSS 1.06402f
C957 a_7399_764.n1 DVSS 3.12204f
C958 a_7399_764.t4 DVSS 1.81038f
C959 a_7399_764.n2 DVSS 0.434584f
C960 a_7399_764.t6 DVSS 1.81038f
C961 a_7399_764.n3 DVSS 0.01455f
C962 a_7399_764.n4 DVSS 3.13034f
C963 a_7399_764.n5 DVSS 1.71545f
C964 a_7399_764.t7 DVSS 1.81038f
C965 a_7399_764.n6 DVSS 0.015267f
C966 a_7399_764.n7 DVSS 1.71363f
C967 a_7399_764.t5 DVSS 1.81038f
C968 a_7399_764.n8 DVSS 1.40668f
C969 a_7399_764.n9 DVSS 0.966925f
C970 a_7399_764.t2 DVSS 9.646111f
C971 a_7399_764.n10 DVSS 0.783271f
C972 a_7399_764.t3 DVSS 1.50783f
C973 a_7399_764.n11 DVSS 1.33404f
C974 a_7399_764.n12 DVSS 0.355312f
C975 a_7399_764.t1 DVSS 0.17422f
C976 a_495_764.t1 DVSS 1.01722f
C977 a_495_764.t2 DVSS 0.819917f
C978 a_495_764.n0 DVSS 7.34093f
C979 a_495_764.t0 DVSS 0.821933f
C980 a_237_764.n0 DVSS 1.10202f
C981 a_237_764.n1 DVSS 0.044802f
C982 a_237_764.n2 DVSS 0.207468f
C983 a_237_764.n3 DVSS 1.47562f
C984 a_237_764.t1 DVSS 0.112149f
C985 a_237_764.t5 DVSS 1.25071f
C986 a_237_764.t6 DVSS 1.25043f
C987 a_237_764.n4 DVSS 0.138379f
C988 a_237_764.t0 DVSS 1.20233f
C989 a_237_764.t2 DVSS 1.20233f
C990 a_237_764.n5 DVSS 0.43999f
C991 a_237_764.n6 DVSS 0.440082f
C992 a_237_764.t4 DVSS 0.992813f
C993 a_237_764.n7 DVSS 0.228721f
C994 a_237_764.t3 DVSS 0.112149f
C995 a_4215_764.t2 DVSS 0.175222f
C996 a_4215_764.n0 DVSS 1.07013f
C997 a_4215_764.n1 DVSS 3.13998f
C998 a_4215_764.t4 DVSS 1.82078f
C999 a_4215_764.n2 DVSS 0.437082f
C1000 a_4215_764.t5 DVSS 1.82078f
C1001 a_4215_764.n3 DVSS 0.014634f
C1002 a_4215_764.n4 DVSS 3.14834f
C1003 a_4215_764.n5 DVSS 1.72531f
C1004 a_4215_764.t6 DVSS 1.82078f
C1005 a_4215_764.n6 DVSS 0.015355f
C1006 a_4215_764.n7 DVSS 1.72348f
C1007 a_4215_764.t7 DVSS 1.82078f
C1008 a_4215_764.n8 DVSS 1.41476f
C1009 a_4215_764.n9 DVSS 0.972482f
C1010 a_4215_764.t1 DVSS 9.70155f
C1011 a_4215_764.n10 DVSS 0.787773f
C1012 a_4215_764.t0 DVSS 1.51649f
C1013 a_4215_764.n11 DVSS 1.34171f
C1014 a_4215_764.n12 DVSS 0.357354f
C1015 a_4215_764.t3 DVSS 0.175222f
C1016 a_3421_764.n0 DVSS 1.09121f
C1017 a_3421_764.n1 DVSS 0.044363f
C1018 a_3421_764.n2 DVSS 0.205434f
C1019 a_3421_764.n3 DVSS 1.46115f
C1020 a_3421_764.t2 DVSS 0.111049f
C1021 a_3421_764.t6 DVSS 1.23845f
C1022 a_3421_764.t5 DVSS 1.23817f
C1023 a_3421_764.n4 DVSS 0.137023f
C1024 a_3421_764.t1 DVSS 1.19055f
C1025 a_3421_764.t3 DVSS 1.19055f
C1026 a_3421_764.n5 DVSS 0.435677f
C1027 a_3421_764.n6 DVSS 0.435767f
C1028 a_3421_764.t0 DVSS 0.98308f
C1029 a_3421_764.n7 DVSS 0.226479f
C1030 a_3421_764.t4 DVSS 0.111049f
C1031 a_10047_764.t1 DVSS 1.30204f
C1032 a_10047_764.t2 DVSS 1.05207f
C1033 a_10047_764.n0 DVSS 9.39639f
C1034 a_10047_764.t0 DVSS 1.04949f
C1035 amp_biases_0.ibias1.n0 DVSS 2.00954f
C1036 amp_biases_0.ibias1.t3 DVSS 0.201678f
C1037 amp_biases_0.ibias1.t2 DVSS 0.201678f
C1038 amp_biases_0.ibias1.n1 DVSS 0.709529f
C1039 amp_biases_0.ibias1.n2 DVSS 1.74963f
C1040 amp_biases_0.ibias1.t5 DVSS 1.7505f
C1041 amp_biases_0.ibias1.n3 DVSS 1.84552f
C1042 amp_biases_0.ibias1.t0 DVSS 1.7505f
C1043 amp_biases_0.ibias1.n4 DVSS 1.43134f
C1044 amp_biases_0.ibias1.t1 DVSS 0.754181f
C1045 amp_biases_0.ibias1.n5 DVSS 2.00078f
C1046 amp_biases_0.ibias1.n6 DVSS 0.472308f
C1047 amp_biases_0.ibias1.t4 DVSS 2.16009f
C1048 amp_biases_0.ibias1.n7 DVSS 5.92716f
C1049 ia_opamp_0.ibias.n0 DVSS 2.39206f
C1050 ia_opamp_0.ibias.n1 DVSS 3.91995f
C1051 ia_opamp_0.ibias.t3 DVSS 0.240068f
C1052 ia_opamp_0.ibias.t2 DVSS 0.240068f
C1053 ia_opamp_0.ibias.n2 DVSS 0.845687f
C1054 ia_opamp_0.ibias.t5 DVSS 2.58003f
C1055 ia_opamp_0.ibias.t4 DVSS 2.08372f
C1056 ia_opamp_0.ibias.n3 DVSS 2.19683f
C1057 ia_opamp_0.ibias.t0 DVSS 2.08372f
C1058 ia_opamp_0.ibias.n4 DVSS 1.70381f
C1059 ia_opamp_0.ibias.t1 DVSS 0.897744f
C1060 ia_opamp_0.ibias.n5 DVSS 2.38286f
C1061 ia_opamp_0.ibias.n6 DVSS 5.30135f
C1062 a_9789_764.n0 DVSS 1.37435f
C1063 a_9789_764.t2 DVSS 0.104452f
C1064 a_9789_764.n1 DVSS 0.155022f
C1065 a_9789_764.t5 DVSS 1.16488f
C1066 a_9789_764.t6 DVSS 1.16462f
C1067 a_9789_764.n2 DVSS 0.128883f
C1068 a_9789_764.n3 DVSS 0.847858f
C1069 a_9789_764.t3 DVSS 1.11982f
C1070 a_9789_764.t1 DVSS 1.11982f
C1071 a_9789_764.n4 DVSS 0.038208f
C1072 a_9789_764.n5 DVSS 0.409795f
C1073 a_9789_764.n6 DVSS 0.409795f
C1074 a_9789_764.n7 DVSS 0.041813f
C1075 a_9789_764.n8 DVSS 0.178532f
C1076 a_9789_764.t0 DVSS 0.924679f
C1077 a_9789_764.n9 DVSS 0.213024f
C1078 a_9789_764.t4 DVSS 0.104452f
C1079 a_204_12823.n0 DVSS 5.21676f
C1080 a_204_12823.n1 DVSS 5.2502f
C1081 a_204_12823.n2 DVSS 8.251611f
C1082 a_204_12823.n3 DVSS 7.84186f
C1083 a_204_12823.n4 DVSS 5.2502f
C1084 a_204_12823.n5 DVSS 0.855365f
C1085 a_204_12823.n6 DVSS 0.187697f
C1086 a_204_12823.t4 DVSS 0.052236f
C1087 a_204_12823.t2 DVSS 0.052236f
C1088 a_204_12823.t3 DVSS 0.314352f
C1089 a_204_12823.t10 DVSS 1.82794f
C1090 a_204_12823.t14 DVSS 1.82794f
C1091 a_204_12823.t13 DVSS 1.82794f
C1092 a_204_12823.t16 DVSS 1.82794f
C1093 a_204_12823.t15 DVSS 1.82794f
C1094 a_204_12823.t6 DVSS 1.83379f
C1095 a_204_12823.t11 DVSS 1.82794f
C1096 a_204_12823.t12 DVSS 1.82794f
C1097 a_204_12823.t5 DVSS 1.82794f
C1098 a_204_12823.t7 DVSS 1.82794f
C1099 a_204_12823.t8 DVSS 1.82794f
C1100 a_204_12823.t9 DVSS 1.83379f
C1101 a_204_12823.t1 DVSS 0.314352f
C1102 a_204_12823.n7 DVSS 0.240629f
C1103 a_204_12823.n8 DVSS 3.94466f
C1104 a_204_12823.t0 DVSS 1.4809f
C1105 a_10583_764.n0 DVSS 4.91904f
C1106 a_10583_764.n1 DVSS 1.08236f
C1107 a_10583_764.n2 DVSS 4.92935f
C1108 a_10583_764.t1 DVSS 0.177224f
C1109 a_10583_764.t4 DVSS 1.84159f
C1110 a_10583_764.n3 DVSS 0.442077f
C1111 a_10583_764.t7 DVSS 1.84159f
C1112 a_10583_764.n4 DVSS 0.014801f
C1113 a_10583_764.t6 DVSS 1.84159f
C1114 a_10583_764.n5 DVSS 0.01553f
C1115 a_10583_764.t5 DVSS 1.84159f
C1116 a_10583_764.n6 DVSS 1.43093f
C1117 a_10583_764.n7 DVSS 0.983596f
C1118 a_10583_764.t2 DVSS 9.81242f
C1119 a_10583_764.n8 DVSS 0.796776f
C1120 a_10583_764.t3 DVSS 1.53383f
C1121 a_10583_764.n9 DVSS 1.35704f
C1122 a_10583_764.n10 DVSS 0.361438f
C1123 a_10583_764.t0 DVSS 0.177224f
C1124 D03v3.t0 DVSS 0.055178f
C1125 D03v3.t3 DVSS 1.23591f
C1126 D03v3.t2 DVSS 1.23945f
C1127 D03v3.n0 DVSS 4.581009f
C1128 D03v3.n1 DVSS 3.85231f
C1129 D03v3.n2 DVSS 0.046538f
C1130 D03v3.t1 DVSS 0.051818f
C1131 D03v3.n3 DVSS 0.045709f
C1132 a_12973_764.n0 DVSS 1.03719f
C1133 a_12973_764.n1 DVSS 0.042167f
C1134 a_12973_764.n2 DVSS 0.195264f
C1135 a_12973_764.n3 DVSS 1.38882f
C1136 a_12973_764.t1 DVSS 0.105552f
C1137 a_12973_764.t5 DVSS 1.17714f
C1138 a_12973_764.t6 DVSS 1.17687f
C1139 a_12973_764.n4 DVSS 0.130239f
C1140 a_12973_764.t2 DVSS 1.13161f
C1141 a_12973_764.t0 DVSS 1.13161f
C1142 a_12973_764.n5 DVSS 0.414109f
C1143 a_12973_764.n6 DVSS 0.414195f
C1144 a_12973_764.t4 DVSS 0.934412f
C1145 a_12973_764.n7 DVSS 0.215267f
C1146 a_12973_764.t3 DVSS 0.105552f
C1147 a_16150_281.t1 DVSS 4.66674f
C1148 a_16150_281.t0 DVSS 0.133257f
C1149 D63v3.n0 DVSS 9.9677f
C1150 D63v3.t0 DVSS 0.043325f
C1151 D63v3.t3 DVSS 1.05171f
C1152 D63v3.n1 DVSS 2.2139f
C1153 D63v3.t5 DVSS 0.984823f
C1154 D63v3.n2 DVSS 1.56275f
C1155 D63v3.t2 DVSS 1.05047f
C1156 D63v3.t4 DVSS 1.04652f
C1157 D63v3.n3 DVSS 0.036541f
C1158 D63v3.t1 DVSS 0.040686f
C1159 D63v3.n4 DVSS 0.03589f
C1160 a_13817_n4916.t10 DVSS 0.229593f
C1161 a_13817_n4916.t7 DVSS 0.051556f
C1162 a_13817_n4916.t8 DVSS 0.051556f
C1163 a_13817_n4916.n0 DVSS 0.148717f
C1164 a_13817_n4916.n1 DVSS 0.548339f
C1165 a_13817_n4916.t5 DVSS 0.051556f
C1166 a_13817_n4916.t12 DVSS 0.051556f
C1167 a_13817_n4916.n2 DVSS 0.148717f
C1168 a_13817_n4916.n3 DVSS 0.292681f
C1169 a_13817_n4916.t9 DVSS 0.051556f
C1170 a_13817_n4916.t13 DVSS 0.051556f
C1171 a_13817_n4916.n4 DVSS 0.148717f
C1172 a_13817_n4916.n5 DVSS 0.389725f
C1173 a_13817_n4916.t11 DVSS 0.180177f
C1174 a_13817_n4916.n6 DVSS 0.473352f
C1175 a_13817_n4916.t2 DVSS 0.082128f
C1176 a_13817_n4916.n7 DVSS 1.35453f
C1177 a_13817_n4916.t4 DVSS 0.082128f
C1178 a_13817_n4916.n8 DVSS 0.802634f
C1179 a_13817_n4916.t1 DVSS 0.082128f
C1180 a_13817_n4916.n9 DVSS 0.802634f
C1181 a_13817_n4916.t14 DVSS 0.082128f
C1182 a_13817_n4916.n10 DVSS 0.802634f
C1183 a_13817_n4916.t3 DVSS 0.082128f
C1184 a_13817_n4916.n11 DVSS 0.802634f
C1185 a_13817_n4916.t6 DVSS 0.082128f
C1186 a_13817_n4916.n12 DVSS 0.802634f
C1187 a_13817_n4916.t15 DVSS 0.082128f
C1188 a_13817_n4916.n13 DVSS 1.20599f
C1189 a_13817_n4916.t0 DVSS 0.382057f
C1190 a_13817_n9984.t6 DVSS 0.227386f
C1191 a_13817_n9984.t11 DVSS 0.051061f
C1192 a_13817_n9984.t9 DVSS 0.051061f
C1193 a_13817_n9984.n0 DVSS 0.147287f
C1194 a_13817_n9984.n1 DVSS 0.543067f
C1195 a_13817_n9984.t5 DVSS 0.051061f
C1196 a_13817_n9984.t7 DVSS 0.051061f
C1197 a_13817_n9984.n2 DVSS 0.147287f
C1198 a_13817_n9984.n3 DVSS 0.289867f
C1199 a_13817_n9984.t10 DVSS 0.051061f
C1200 a_13817_n9984.t13 DVSS 0.051061f
C1201 a_13817_n9984.n4 DVSS 0.147287f
C1202 a_13817_n9984.n5 DVSS 0.385977f
C1203 a_13817_n9984.t12 DVSS 0.178445f
C1204 a_13817_n9984.n6 DVSS 0.4688f
C1205 a_13817_n9984.t15 DVSS 0.081338f
C1206 a_13817_n9984.n7 DVSS 1.3415f
C1207 a_13817_n9984.t1 DVSS 0.081338f
C1208 a_13817_n9984.n8 DVSS 0.794916f
C1209 a_13817_n9984.t3 DVSS 0.081338f
C1210 a_13817_n9984.n9 DVSS 0.794916f
C1211 a_13817_n9984.t14 DVSS 0.081338f
C1212 a_13817_n9984.n10 DVSS 0.794916f
C1213 a_13817_n9984.t2 DVSS 0.081338f
C1214 a_13817_n9984.n11 DVSS 0.794916f
C1215 a_13817_n9984.t8 DVSS 0.081338f
C1216 a_13817_n9984.n12 DVSS 0.794916f
C1217 a_13817_n9984.t4 DVSS 0.081338f
C1218 a_13817_n9984.n13 DVSS 1.1944f
C1219 a_13817_n9984.t0 DVSS 0.378383f
C1220 a_6605_764.n0 DVSS 1.02639f
C1221 a_6605_764.n1 DVSS 0.041727f
C1222 a_6605_764.n2 DVSS 0.19323f
C1223 a_6605_764.n3 DVSS 1.37435f
C1224 a_6605_764.t1 DVSS 0.104452f
C1225 a_6605_764.t5 DVSS 1.16488f
C1226 a_6605_764.t6 DVSS 1.16462f
C1227 a_6605_764.n4 DVSS 0.128883f
C1228 a_6605_764.t2 DVSS 1.11982f
C1229 a_6605_764.t0 DVSS 1.11982f
C1230 a_6605_764.n5 DVSS 0.409795f
C1231 a_6605_764.n6 DVSS 0.40988f
C1232 a_6605_764.t4 DVSS 0.924679f
C1233 a_6605_764.n7 DVSS 0.213024f
C1234 a_6605_764.t3 DVSS 0.104452f
C1235 a_16157_764.n0 DVSS 1.01559f
C1236 a_16157_764.n1 DVSS 0.041288f
C1237 a_16157_764.n2 DVSS 0.191196f
C1238 a_16157_764.n3 DVSS 1.35989f
C1239 a_16157_764.t1 DVSS 0.103353f
C1240 a_16157_764.t6 DVSS 1.15262f
C1241 a_16157_764.t5 DVSS 1.15236f
C1242 a_16157_764.n4 DVSS 0.127526f
C1243 a_16157_764.t0 DVSS 1.10803f
C1244 a_16157_764.t2 DVSS 1.10803f
C1245 a_16157_764.n5 DVSS 0.405481f
C1246 a_16157_764.n6 DVSS 0.405566f
C1247 a_16157_764.t4 DVSS 0.914945f
C1248 a_16157_764.n7 DVSS 0.210782f
C1249 a_16157_764.t3 DVSS 0.103353f
C1250 a_230_281.t1 DVSS 4.66674f
C1251 a_230_281.t0 DVSS 0.133257f
C1252 a_12405_n4916.t6 DVSS 0.206656f
C1253 a_12405_n4916.t4 DVSS 0.045806f
C1254 a_12405_n4916.t5 DVSS 0.045806f
C1255 a_12405_n4916.n0 DVSS 0.133456f
C1256 a_12405_n4916.n1 DVSS 0.55826f
C1257 a_12405_n4916.t3 DVSS 0.161009f
C1258 a_12405_n4916.n2 DVSS 0.38851f
C1259 a_12405_n4916.t1 DVSS 0.068731f
C1260 a_12405_n4916.n3 DVSS 1.0536f
C1261 a_12405_n4916.t2 DVSS 0.068731f
C1262 a_12405_n4916.n4 DVSS 0.671705f
C1263 a_12405_n4916.t7 DVSS 0.068731f
C1264 a_12405_n4916.n5 DVSS 1.00927f
C1265 a_12405_n4916.t0 DVSS 0.319734f
C1266 x8.V2.t70 DVSS 1.02048f
C1267 x8.V2.t45 DVSS 0.10721f
C1268 x8.V2.t35 DVSS 0.10721f
C1269 x8.V2.n0 DVSS 0.21866f
C1270 x8.V2.n1 DVSS 0.431955f
C1271 x8.V2.n2 DVSS 0.134909f
C1272 x8.V2.n3 DVSS 0.19669f
C1273 x8.V2.t62 DVSS 0.032192f
C1274 x8.V2.n4 DVSS 0.280494f
C1275 x8.V2.t17 DVSS 0.032192f
C1276 x8.V2.n5 DVSS 0.19669f
C1277 x8.V2.t23 DVSS 0.032192f
C1278 x8.V2.n6 DVSS 0.280494f
C1279 x8.V2.t50 DVSS 0.032192f
C1280 x8.V2.n7 DVSS 0.19669f
C1281 x8.V2.t2 DVSS 0.032192f
C1282 x8.V2.n8 DVSS 0.280494f
C1283 x8.V2.t9 DVSS 0.032192f
C1284 x8.V2.n9 DVSS 0.19669f
C1285 x8.V2.t10 DVSS 0.032192f
C1286 x8.V2.n10 DVSS 0.280494f
C1287 x8.V2.t12 DVSS 0.032192f
C1288 x8.V2.n11 DVSS 0.19669f
C1289 x8.V2.t44 DVSS 0.032192f
C1290 x8.V2.n12 DVSS 0.280494f
C1291 x8.V2.t55 DVSS 0.032192f
C1292 x8.V2.n13 DVSS 0.19669f
C1293 x8.V2.t24 DVSS 0.032192f
C1294 x8.V2.n14 DVSS 0.280494f
C1295 x8.V2.t13 DVSS 0.032192f
C1296 x8.V2.t20 DVSS 0.169761f
C1297 x8.V2.t33 DVSS 0.115997f
C1298 x8.V2.n15 DVSS 0.105949f
C1299 x8.V2.t59 DVSS 0.115997f
C1300 x8.V2.n16 DVSS 0.10003f
C1301 x8.V2.t31 DVSS 0.115997f
C1302 x8.V2.n17 DVSS 0.10003f
C1303 x8.V2.t26 DVSS 0.032192f
C1304 x8.V2.n18 DVSS 0.285046f
C1305 x8.V2.n19 DVSS 0.116508f
C1306 x8.V2.n20 DVSS 0.328974f
C1307 x8.V2.n21 DVSS 0.280494f
C1308 x8.V2.t36 DVSS 0.032192f
C1309 x8.V2.n22 DVSS 0.280494f
C1310 x8.V2.t0 DVSS 0.115997f
C1311 x8.V2.n23 DVSS 0.19669f
C1312 x8.V2.n24 DVSS 0.19669f
C1313 x8.V2.n25 DVSS 0.19669f
C1314 x8.V2.n26 DVSS 0.19669f
C1315 x8.V2.n27 DVSS 0.280494f
C1316 x8.V2.t67 DVSS 0.032192f
C1317 x8.V2.n28 DVSS 0.280494f
C1318 x8.V2.t60 DVSS 0.032192f
C1319 x8.V2.n29 DVSS 0.280494f
C1320 x8.V2.n30 DVSS 0.19669f
C1321 x8.V2.n31 DVSS 0.19669f
C1322 x8.V2.n32 DVSS 0.19669f
C1323 x8.V2.n33 DVSS 0.280494f
C1324 x8.V2.t49 DVSS 0.032192f
C1325 x8.V2.n34 DVSS 0.280494f
C1326 x8.V2.t25 DVSS 0.032192f
C1327 x8.V2.n35 DVSS 0.280494f
C1328 x8.V2.n36 DVSS 0.19669f
C1329 x8.V2.n37 DVSS 0.19669f
C1330 x8.V2.n38 DVSS 0.19669f
C1331 x8.V2.n39 DVSS 0.280494f
C1332 x8.V2.t56 DVSS 0.032192f
C1333 x8.V2.n40 DVSS 0.280494f
C1334 x8.V2.t29 DVSS 0.032192f
C1335 x8.V2.n41 DVSS 0.280494f
C1336 x8.V2.n42 DVSS 0.19669f
C1337 x8.V2.n43 DVSS 0.19669f
C1338 x8.V2.n44 DVSS 0.19669f
C1339 x8.V2.n45 DVSS 0.280494f
C1340 x8.V2.t3 DVSS 0.032192f
C1341 x8.V2.n46 DVSS 0.280494f
C1342 x8.V2.t52 DVSS 0.032192f
C1343 x8.V2.n47 DVSS 0.280494f
C1344 x8.V2.n48 DVSS 0.19669f
C1345 x8.V2.n49 DVSS 0.19669f
C1346 x8.V2.n50 DVSS 0.19669f
C1347 x8.V2.n51 DVSS 0.280494f
C1348 x8.V2.t41 DVSS 0.032192f
C1349 x8.V2.n52 DVSS 0.280494f
C1350 x8.V2.t63 DVSS 0.032192f
C1351 x8.V2.t40 DVSS 0.032192f
C1352 x8.V2.t11 DVSS 0.032192f
C1353 x8.V2.t21 DVSS 0.032192f
C1354 x8.V2.n53 DVSS 0.280494f
C1355 x8.V2.n54 DVSS 0.19669f
C1356 x8.V2.t43 DVSS 0.032192f
C1357 x8.V2.t5 DVSS 0.032192f
C1358 x8.V2.t65 DVSS 0.032192f
C1359 x8.V2.t38 DVSS 0.032192f
C1360 x8.V2.n55 DVSS 0.280494f
C1361 x8.V2.n56 DVSS 0.19669f
C1362 x8.V2.t7 DVSS 0.032192f
C1363 x8.V2.t58 DVSS 0.032192f
C1364 x8.V2.t6 DVSS 0.032192f
C1365 x8.V2.t57 DVSS 0.032192f
C1366 x8.V2.n57 DVSS 0.280494f
C1367 x8.V2.n58 DVSS 0.19669f
C1368 x8.V2.t47 DVSS 0.032192f
C1369 x8.V2.t66 DVSS 0.032192f
C1370 x8.V2.t39 DVSS 0.032192f
C1371 x8.V2.t68 DVSS 0.032192f
C1372 x8.V2.n59 DVSS 0.280494f
C1373 x8.V2.n60 DVSS 0.19669f
C1374 x8.V2.t1 DVSS 0.032192f
C1375 x8.V2.t19 DVSS 0.032192f
C1376 x8.V2.t54 DVSS 0.032192f
C1377 x8.V2.t28 DVSS 0.032192f
C1378 x8.V2.n61 DVSS 0.280494f
C1379 x8.V2.n62 DVSS 0.19669f
C1380 x8.V2.t15 DVSS 0.032192f
C1381 x8.V2.t64 DVSS 0.032192f
C1382 x8.V2.t61 DVSS 0.032192f
C1383 x8.V2.t14 DVSS 0.032192f
C1384 x8.V2.n63 DVSS 0.280494f
C1385 x8.V2.n64 DVSS 0.19669f
C1386 x8.V2.t4 DVSS 0.032192f
C1387 x8.V2.t27 DVSS 0.032192f
C1388 x8.V2.t22 DVSS 0.032192f
C1389 x8.V2.t18 DVSS 0.032192f
C1390 x8.V2.n65 DVSS 0.280494f
C1391 x8.V2.n66 DVSS 0.19669f
C1392 x8.V2.t37 DVSS 0.032192f
C1393 x8.V2.t51 DVSS 0.032192f
C1394 x8.V2.t16 DVSS 0.032192f
C1395 x8.V2.t8 DVSS 0.032192f
C1396 x8.V2.n67 DVSS 0.280494f
C1397 x8.V2.n68 DVSS 0.378131f
C1398 x8.V2.t69 DVSS 0.032192f
C1399 x8.V2.t42 DVSS 0.032192f
C1400 x8.V2.t48 DVSS 0.032192f
C1401 x8.V2.t53 DVSS 0.040211f
C1402 x8.V2.n69 DVSS 0.40372f
C1403 x8.V2.n70 DVSS 0.280494f
C1404 x8.V2.n71 DVSS 0.280494f
C1405 x8.V2.n72 DVSS 0.280494f
C1406 x8.V2.n73 DVSS 0.19669f
C1407 x8.V2.n74 DVSS 0.19669f
C1408 x8.V2.n75 DVSS 0.19669f
C1409 x8.V2.n76 DVSS 0.280494f
C1410 x8.V2.n77 DVSS 0.280494f
C1411 x8.V2.n78 DVSS 0.280494f
C1412 x8.V2.n79 DVSS 0.19669f
C1413 x8.V2.n80 DVSS 0.19669f
C1414 x8.V2.n81 DVSS 0.19669f
C1415 x8.V2.n82 DVSS 0.280494f
C1416 x8.V2.n83 DVSS 0.280494f
C1417 x8.V2.n84 DVSS 0.280494f
C1418 x8.V2.n85 DVSS 0.19669f
C1419 x8.V2.n86 DVSS 0.19669f
C1420 x8.V2.n87 DVSS 0.19669f
C1421 x8.V2.n88 DVSS 0.280494f
C1422 x8.V2.n89 DVSS 0.280494f
C1423 x8.V2.n90 DVSS 0.280494f
C1424 x8.V2.n91 DVSS 0.19669f
C1425 x8.V2.n92 DVSS 0.19669f
C1426 x8.V2.n93 DVSS 0.19669f
C1427 x8.V2.n94 DVSS 0.280494f
C1428 x8.V2.n95 DVSS 0.280494f
C1429 x8.V2.n96 DVSS 0.280494f
C1430 x8.V2.n97 DVSS 0.19669f
C1431 x8.V2.n98 DVSS 0.19669f
C1432 x8.V2.n99 DVSS 0.19669f
C1433 x8.V2.n100 DVSS 0.280494f
C1434 x8.V2.n101 DVSS 0.280494f
C1435 x8.V2.n102 DVSS 0.280494f
C1436 x8.V2.n103 DVSS 0.19669f
C1437 x8.V2.n104 DVSS 0.19669f
C1438 x8.V2.n105 DVSS 0.19669f
C1439 x8.V2.n106 DVSS 0.280494f
C1440 x8.V2.n107 DVSS 0.280494f
C1441 x8.V2.n108 DVSS 0.280494f
C1442 x8.V2.n109 DVSS 0.19669f
C1443 x8.V2.n110 DVSS 0.19669f
C1444 x8.V2.n111 DVSS 0.19669f
C1445 x8.V2.n112 DVSS 0.280494f
C1446 x8.V2.n113 DVSS 0.280494f
C1447 x8.V2.n114 DVSS 0.280494f
C1448 x8.V2.n115 DVSS 0.19669f
C1449 x8.V2.n116 DVSS 0.19669f
C1450 x8.V2.n117 DVSS 0.19669f
C1451 x8.V2.n118 DVSS 0.280494f
C1452 x8.V2.n119 DVSS 0.280494f
C1453 x8.V2.n120 DVSS 0.280494f
C1454 x8.V2.n121 DVSS 0.160126f
C1455 x8.V2.n122 DVSS 1.40541f
C1456 x8.V2.n123 DVSS 1.83456f
C1457 x8.V2.t34 DVSS 0.10721f
C1458 x8.V2.t46 DVSS 0.10721f
C1459 x8.V2.n124 DVSS 0.21866f
C1460 x8.V2.n125 DVSS 0.417768f
C1461 x8.V2.n126 DVSS 0.443311f
C1462 x8.V2.n127 DVSS 0.158637f
C1463 x8.V2.t32 DVSS 0.226759f
C1464 x8.V2.t30 DVSS 0.3749f
C1465 x8.V2.n128 DVSS 0.849774f
C1466 x8.V2.n129 DVSS 0.875421f
C1467 x8.V2.n130 DVSS 0.473817f
C1468 a_3720_n4916.t9 DVSS 0.21414f
C1469 a_3720_n4916.t6 DVSS 0.048086f
C1470 a_3720_n4916.t5 DVSS 0.048086f
C1471 a_3720_n4916.n0 DVSS 0.138707f
C1472 a_3720_n4916.n1 DVSS 0.511432f
C1473 a_3720_n4916.t3 DVSS 0.048086f
C1474 a_3720_n4916.t4 DVSS 0.048086f
C1475 a_3720_n4916.n2 DVSS 0.138707f
C1476 a_3720_n4916.n3 DVSS 0.272982f
C1477 a_3720_n4916.t7 DVSS 0.048086f
C1478 a_3720_n4916.t2 DVSS 0.048086f
C1479 a_3720_n4916.n4 DVSS 0.138707f
C1480 a_3720_n4916.n5 DVSS 0.363493f
C1481 a_3720_n4916.t8 DVSS 0.16805f
C1482 a_3720_n4916.n6 DVSS 0.441492f
C1483 a_3720_n4916.t10 DVSS 0.0766f
C1484 a_3720_n4916.n7 DVSS 1.26336f
C1485 a_3720_n4916.t15 DVSS 0.0766f
C1486 a_3720_n4916.n8 DVSS 0.748611f
C1487 a_3720_n4916.t13 DVSS 0.0766f
C1488 a_3720_n4916.n9 DVSS 0.748611f
C1489 a_3720_n4916.t12 DVSS 0.0766f
C1490 a_3720_n4916.n10 DVSS 0.748611f
C1491 a_3720_n4916.t11 DVSS 0.0766f
C1492 a_3720_n4916.n11 DVSS 0.748611f
C1493 a_3720_n4916.t1 DVSS 0.0766f
C1494 a_3720_n4916.n12 DVSS 0.748611f
C1495 a_3720_n4916.t14 DVSS 0.0766f
C1496 a_3720_n4916.n13 DVSS 1.12482f
C1497 a_3720_n4916.t0 DVSS 0.356341f
C1498 a_12405_n9984.t5 DVSS 0.223877f
C1499 a_12405_n9984.t3 DVSS 0.049623f
C1500 a_12405_n9984.t4 DVSS 0.049623f
C1501 a_12405_n9984.n0 DVSS 0.144577f
C1502 a_12405_n9984.n1 DVSS 0.604781f
C1503 a_12405_n9984.t2 DVSS 0.174426f
C1504 a_12405_n9984.n2 DVSS 0.420886f
C1505 a_12405_n9984.t1 DVSS 0.074458f
C1506 a_12405_n9984.n3 DVSS 1.1414f
C1507 a_12405_n9984.t6 DVSS 0.076501f
C1508 a_12405_n9984.t7 DVSS 0.074458f
C1509 a_12405_n9984.n4 DVSS 1.36325f
C1510 a_12405_n9984.n5 DVSS 0.472237f
C1511 a_12405_n9984.t0 DVSS 0.329902f
C1512 D73v3.n0 DVSS 6.15118f
C1513 D73v3.n1 DVSS 8.740789f
C1514 D73v3.t0 DVSS 0.049266f
C1515 D73v3.t3 DVSS 1.08453f
C1516 D73v3.t9 DVSS 1.15894f
C1517 D73v3.t7 DVSS 1.15303f
C1518 D73v3.t5 DVSS 1.15299f
C1519 D73v3.n2 DVSS 1.76094f
C1520 D73v3.t8 DVSS 1.15894f
C1521 D73v3.t6 DVSS 1.15303f
C1522 D73v3.t4 DVSS 1.15299f
C1523 D73v3.t2 DVSS 1.15299f
C1524 D73v3.n3 DVSS 6.48345f
C1525 D73v3.n4 DVSS 0.041552f
C1526 D73v3.t1 DVSS 0.046266f
C1527 D73v3.n5 DVSS 0.040812f
C1528 AVOUT1.t6 DVSS 0.168733f
C1529 AVOUT1.t7 DVSS 0.168733f
C1530 AVOUT1.n0 DVSS 0.542636f
C1531 AVOUT1.t12 DVSS 0.168733f
C1532 AVOUT1.t13 DVSS 0.168733f
C1533 AVOUT1.n1 DVSS 0.535748f
C1534 AVOUT1.n2 DVSS 1.55776f
C1535 AVOUT1.t38 DVSS 1.60594f
C1536 AVOUT1.n3 DVSS 1.63804f
C1537 AVOUT1.t22 DVSS 0.061837f
C1538 AVOUT1.n4 DVSS 1.48554f
C1539 AVOUT1.t0 DVSS 0.061837f
C1540 AVOUT1.n5 DVSS 0.604967f
C1541 AVOUT1.t32 DVSS 0.061837f
C1542 AVOUT1.n6 DVSS 0.604967f
C1543 AVOUT1.t25 DVSS 0.061837f
C1544 AVOUT1.n7 DVSS 0.604967f
C1545 AVOUT1.t28 DVSS 0.061837f
C1546 AVOUT1.n8 DVSS 0.604967f
C1547 AVOUT1.t21 DVSS 0.061837f
C1548 AVOUT1.n9 DVSS 0.604967f
C1549 AVOUT1.t18 DVSS 0.061837f
C1550 AVOUT1.n10 DVSS 0.604967f
C1551 AVOUT1.t26 DVSS 0.061837f
C1552 AVOUT1.n11 DVSS 0.604967f
C1553 AVOUT1.t8 DVSS 0.061837f
C1554 AVOUT1.n12 DVSS 0.604967f
C1555 AVOUT1.t1 DVSS 0.061837f
C1556 AVOUT1.n13 DVSS 0.604967f
C1557 AVOUT1.t29 DVSS 0.061837f
C1558 AVOUT1.n14 DVSS 0.604967f
C1559 AVOUT1.t4 DVSS 0.061837f
C1560 AVOUT1.n15 DVSS 0.604967f
C1561 AVOUT1.t2 DVSS 0.061837f
C1562 AVOUT1.n16 DVSS 0.604967f
C1563 AVOUT1.t17 DVSS 0.061837f
C1564 AVOUT1.n17 DVSS 0.604967f
C1565 AVOUT1.t33 DVSS 0.061837f
C1566 AVOUT1.n18 DVSS 0.585628f
C1567 AVOUT1.n19 DVSS 0.273693f
C1568 AVOUT1.t11 DVSS 0.062137f
C1569 AVOUT1.n20 DVSS 0.566774f
C1570 AVOUT1.t35 DVSS 0.061837f
C1571 AVOUT1.n21 DVSS 0.748071f
C1572 AVOUT1.t15 DVSS 0.061837f
C1573 AVOUT1.n22 DVSS 0.879573f
C1574 AVOUT1.t34 DVSS 0.061837f
C1575 AVOUT1.n23 DVSS 0.604967f
C1576 AVOUT1.t20 DVSS 0.061837f
C1577 AVOUT1.n24 DVSS 0.604967f
C1578 AVOUT1.t19 DVSS 0.061837f
C1579 AVOUT1.n25 DVSS 0.501828f
C1580 AVOUT1.n26 DVSS 0.307968f
C1581 AVOUT1.t16 DVSS 0.061837f
C1582 AVOUT1.n27 DVSS 0.557265f
C1583 AVOUT1.t9 DVSS 0.061837f
C1584 AVOUT1.n28 DVSS 0.604967f
C1585 AVOUT1.t24 DVSS 0.061837f
C1586 AVOUT1.n29 DVSS 0.604967f
C1587 AVOUT1.t3 DVSS 0.061837f
C1588 AVOUT1.n30 DVSS 0.938877f
C1589 AVOUT1.t10 DVSS 0.061837f
C1590 AVOUT1.n31 DVSS 0.938877f
C1591 AVOUT1.t36 DVSS 0.061837f
C1592 AVOUT1.n32 DVSS 0.604967f
C1593 AVOUT1.t14 DVSS 0.061837f
C1594 AVOUT1.n33 DVSS 0.604967f
C1595 AVOUT1.t31 DVSS 0.061837f
C1596 AVOUT1.n34 DVSS 0.9002f
C1597 AVOUT1.t37 DVSS 0.061837f
C1598 AVOUT1.n35 DVSS 0.9002f
C1599 AVOUT1.t5 DVSS 0.061837f
C1600 AVOUT1.n36 DVSS 0.861523f
C1601 AVOUT1.t30 DVSS 0.061837f
C1602 AVOUT1.n37 DVSS 1.05104f
C1603 AVOUT1.t23 DVSS 0.061837f
C1604 AVOUT1.n38 DVSS 0.765579f
C1605 AVOUT1.n39 DVSS 0.055549f
C1606 AVOUT1.n40 DVSS 0.74356f
C1607 AVOUT1.n41 DVSS 1.2835f
C1608 AVOUT1.n42 DVSS 0.782372f
C1609 AVOUT1.t27 DVSS 0.59004f
C1610 AVOUT1.n43 DVSS 1.63395f
C1611 AVOUT1.n44 DVSS 1.68859f
C1612 a_6164_n4916.t11 DVSS 0.211333f
C1613 a_6164_n4916.t5 DVSS 0.047738f
C1614 a_6164_n4916.t12 DVSS 0.047738f
C1615 a_6164_n4916.n0 DVSS 0.137856f
C1616 a_6164_n4916.n1 DVSS 0.495309f
C1617 a_6164_n4916.t17 DVSS 0.047738f
C1618 a_6164_n4916.t6 DVSS 0.047738f
C1619 a_6164_n4916.n2 DVSS 0.137856f
C1620 a_6164_n4916.n3 DVSS 0.270326f
C1621 a_6164_n4916.t14 DVSS 0.047738f
C1622 a_6164_n4916.t13 DVSS 0.047738f
C1623 a_6164_n4916.n4 DVSS 0.137856f
C1624 a_6164_n4916.n5 DVSS 0.270326f
C1625 a_6164_n4916.t8 DVSS 0.047738f
C1626 a_6164_n4916.t7 DVSS 0.047738f
C1627 a_6164_n4916.n6 DVSS 0.137856f
C1628 a_6164_n4916.n7 DVSS 0.270326f
C1629 a_6164_n4916.t15 DVSS 0.047738f
C1630 a_6164_n4916.t18 DVSS 0.047738f
C1631 a_6164_n4916.n8 DVSS 0.137856f
C1632 a_6164_n4916.n9 DVSS 0.270476f
C1633 a_6164_n4916.t9 DVSS 0.047738f
C1634 a_6164_n4916.t16 DVSS 0.047738f
C1635 a_6164_n4916.n10 DVSS 0.137856f
C1636 a_6164_n4916.n11 DVSS 0.360307f
C1637 a_6164_n4916.t10 DVSS 0.166942f
C1638 a_6164_n4916.n12 DVSS 0.504931f
C1639 a_6164_n4916.t22 DVSS 0.0757f
C1640 a_6164_n4916.n13 DVSS 1.04845f
C1641 a_6164_n4916.t29 DVSS 0.077778f
C1642 a_6164_n4916.t28 DVSS 0.0757f
C1643 a_6164_n4916.n14 DVSS 1.38909f
C1644 a_6164_n4916.t19 DVSS 0.0757f
C1645 a_6164_n4916.n15 DVSS 0.740686f
C1646 a_6164_n4916.t2 DVSS 0.0757f
C1647 a_6164_n4916.n16 DVSS 0.740686f
C1648 a_6164_n4916.t3 DVSS 0.0757f
C1649 a_6164_n4916.n17 DVSS 0.740686f
C1650 a_6164_n4916.t26 DVSS 0.0757f
C1651 a_6164_n4916.n18 DVSS 0.740686f
C1652 a_6164_n4916.t1 DVSS 0.0757f
C1653 a_6164_n4916.n19 DVSS 0.740686f
C1654 a_6164_n4916.t4 DVSS 0.0757f
C1655 a_6164_n4916.n20 DVSS 0.740686f
C1656 a_6164_n4916.t24 DVSS 0.0757f
C1657 a_6164_n4916.n21 DVSS 0.740686f
C1658 a_6164_n4916.t20 DVSS 0.0757f
C1659 a_6164_n4916.n22 DVSS 0.740686f
C1660 a_6164_n4916.t21 DVSS 0.0757f
C1661 a_6164_n4916.n23 DVSS 0.740686f
C1662 a_6164_n4916.t25 DVSS 0.0757f
C1663 a_6164_n4916.n24 DVSS 0.740686f
C1664 a_6164_n4916.t23 DVSS 0.0757f
C1665 a_6164_n4916.n25 DVSS 0.740686f
C1666 a_6164_n4916.t27 DVSS 0.0757f
C1667 a_6164_n4916.n26 DVSS 0.740686f
C1668 a_6164_n4916.n27 DVSS 0.480985f
C1669 a_6164_n4916.t0 DVSS 0.335401f
C1670 a_3720_n9984.t10 DVSS 0.231801f
C1671 a_3720_n9984.t7 DVSS 0.052052f
C1672 a_3720_n9984.t6 DVSS 0.052052f
C1673 a_3720_n9984.n0 DVSS 0.150147f
C1674 a_3720_n9984.n1 DVSS 0.553612f
C1675 a_3720_n9984.t4 DVSS 0.052052f
C1676 a_3720_n9984.t5 DVSS 0.052052f
C1677 a_3720_n9984.n2 DVSS 0.150147f
C1678 a_3720_n9984.n3 DVSS 0.295496f
C1679 a_3720_n9984.t8 DVSS 0.052052f
C1680 a_3720_n9984.t3 DVSS 0.052052f
C1681 a_3720_n9984.n4 DVSS 0.150147f
C1682 a_3720_n9984.n5 DVSS 0.393472f
C1683 a_3720_n9984.t9 DVSS 0.18191f
C1684 a_3720_n9984.n6 DVSS 0.477903f
C1685 a_3720_n9984.t11 DVSS 0.082918f
C1686 a_3720_n9984.n7 DVSS 1.36755f
C1687 a_3720_n9984.t12 DVSS 0.082918f
C1688 a_3720_n9984.n8 DVSS 0.810352f
C1689 a_3720_n9984.t15 DVSS 0.082918f
C1690 a_3720_n9984.n9 DVSS 0.810352f
C1691 a_3720_n9984.t13 DVSS 0.082918f
C1692 a_3720_n9984.n10 DVSS 0.810352f
C1693 a_3720_n9984.t2 DVSS 0.082918f
C1694 a_3720_n9984.n11 DVSS 0.810352f
C1695 a_3720_n9984.t1 DVSS 0.082918f
C1696 a_3720_n9984.n12 DVSS 0.810352f
C1697 a_3720_n9984.t14 DVSS 0.085192f
C1698 a_3720_n9984.n13 DVSS 1.23366f
C1699 a_3720_n9984.t0 DVSS 0.367381f
C1700 D33v3.n0 DVSS 11.9137f
C1701 D33v3.n1 DVSS 11.4176f
C1702 D33v3.t0 DVSS 0.044682f
C1703 D33v3.t5 DVSS 1.01167f
C1704 D33v3.t7 DVSS 1.00631f
C1705 D33v3.t17 DVSS 1.00631f
C1706 D33v3.t15 DVSS 1.00631f
C1707 D33v3.t13 DVSS 1.00631f
C1708 D33v3.t9 DVSS 1.00631f
C1709 D33v3.t11 DVSS 1.00631f
C1710 D33v3.t3 DVSS 0.944057f
C1711 D33v3.t2 DVSS 0.944894f
C1712 D33v3.t4 DVSS 1.01167f
C1713 D33v3.t6 DVSS 1.00631f
C1714 D33v3.t16 DVSS 1.00631f
C1715 D33v3.t14 DVSS 1.00631f
C1716 D33v3.t12 DVSS 1.00631f
C1717 D33v3.t8 DVSS 1.00631f
C1718 D33v3.t10 DVSS 1.00631f
C1719 D33v3.n2 DVSS 3.28353f
C1720 D33v3.n3 DVSS 3.083f
C1721 D33v3.n4 DVSS 0.037686f
C1722 D33v3.t1 DVSS 0.041961f
C1723 D33v3.n5 DVSS 0.037014f
C1724 AVOUT2.t38 DVSS 1.44051f
C1725 AVOUT2.n0 DVSS 2.02366f
C1726 AVOUT2.t27 DVSS 0.150038f
C1727 AVOUT2.t5 DVSS 0.151352f
C1728 AVOUT2.t24 DVSS 0.151352f
C1729 AVOUT2.n1 DVSS 0.486739f
C1730 AVOUT2.t23 DVSS 0.151352f
C1731 AVOUT2.t4 DVSS 0.151352f
C1732 AVOUT2.n2 DVSS 0.480561f
C1733 AVOUT2.n3 DVSS 1.39729f
C1734 AVOUT2.n4 DVSS 1.5138f
C1735 AVOUT2.t6 DVSS 0.52926f
C1736 AVOUT2.n5 DVSS 1.67475f
C1737 AVOUT2.n6 DVSS 0.952463f
C1738 AVOUT2.n7 DVSS 3.84681f
C1739 AVOUT2.t32 DVSS 0.057f
C1740 AVOUT2.t17 DVSS 0.055467f
C1741 AVOUT2.n8 DVSS 1.01669f
C1742 AVOUT2.t29 DVSS 0.055467f
C1743 AVOUT2.n9 DVSS 0.54265f
C1744 AVOUT2.t3 DVSS 0.055467f
C1745 AVOUT2.n10 DVSS 0.54265f
C1746 AVOUT2.t10 DVSS 0.055467f
C1747 AVOUT2.n11 DVSS 0.54265f
C1748 AVOUT2.t9 DVSS 0.055467f
C1749 AVOUT2.n12 DVSS 0.54265f
C1750 AVOUT2.t12 DVSS 0.055467f
C1751 AVOUT2.n13 DVSS 0.54265f
C1752 AVOUT2.t20 DVSS 0.055467f
C1753 AVOUT2.n14 DVSS 0.54265f
C1754 AVOUT2.t13 DVSS 0.055467f
C1755 AVOUT2.n15 DVSS 0.54265f
C1756 AVOUT2.t26 DVSS 0.055467f
C1757 AVOUT2.n16 DVSS 0.54265f
C1758 AVOUT2.t35 DVSS 0.055467f
C1759 AVOUT2.n17 DVSS 0.54265f
C1760 AVOUT2.t33 DVSS 0.055467f
C1761 AVOUT2.n18 DVSS 0.54265f
C1762 AVOUT2.t18 DVSS 0.055467f
C1763 AVOUT2.n19 DVSS 0.54265f
C1764 AVOUT2.t0 DVSS 0.055467f
C1765 AVOUT2.n20 DVSS 0.54265f
C1766 AVOUT2.t31 DVSS 0.055467f
C1767 AVOUT2.n21 DVSS 0.54265f
C1768 AVOUT2.t25 DVSS 0.055467f
C1769 AVOUT2.n22 DVSS 0.520098f
C1770 AVOUT2.n23 DVSS 2.08182f
C1771 AVOUT2.t16 DVSS 0.055467f
C1772 AVOUT2.n24 DVSS 0.676215f
C1773 AVOUT2.t21 DVSS 0.055467f
C1774 AVOUT2.n25 DVSS 0.54265f
C1775 AVOUT2.t36 DVSS 0.055467f
C1776 AVOUT2.n26 DVSS 0.54265f
C1777 AVOUT2.t22 DVSS 0.055467f
C1778 AVOUT2.n27 DVSS 0.54265f
C1779 AVOUT2.t8 DVSS 0.055467f
C1780 AVOUT2.n28 DVSS 0.54265f
C1781 AVOUT2.t2 DVSS 0.055467f
C1782 AVOUT2.n29 DVSS 0.54265f
C1783 AVOUT2.t1 DVSS 0.055467f
C1784 AVOUT2.n30 DVSS 0.54265f
C1785 AVOUT2.t34 DVSS 0.055467f
C1786 AVOUT2.n31 DVSS 0.842164f
C1787 AVOUT2.t7 DVSS 0.055467f
C1788 AVOUT2.n32 DVSS 0.842164f
C1789 AVOUT2.t14 DVSS 0.055467f
C1790 AVOUT2.n33 DVSS 0.54265f
C1791 AVOUT2.t37 DVSS 0.055467f
C1792 AVOUT2.n34 DVSS 0.54265f
C1793 AVOUT2.t28 DVSS 0.055467f
C1794 AVOUT2.n35 DVSS 0.807471f
C1795 AVOUT2.t30 DVSS 0.055467f
C1796 AVOUT2.n36 DVSS 0.807471f
C1797 AVOUT2.t11 DVSS 0.055467f
C1798 AVOUT2.n37 DVSS 0.772778f
C1799 AVOUT2.t19 DVSS 0.055467f
C1800 AVOUT2.n38 DVSS 0.942773f
C1801 AVOUT2.t15 DVSS 0.055467f
C1802 AVOUT2.n39 DVSS 0.686718f
C1803 AVOUT2.n40 DVSS 0.056839f
C1804 a_6164_n9984.t10 DVSS 0.217371f
C1805 a_6164_n9984.t4 DVSS 0.049102f
C1806 a_6164_n9984.t11 DVSS 0.049102f
C1807 a_6164_n9984.n0 DVSS 0.141794f
C1808 a_6164_n9984.n1 DVSS 0.509461f
C1809 a_6164_n9984.t16 DVSS 0.049102f
C1810 a_6164_n9984.t5 DVSS 0.049102f
C1811 a_6164_n9984.n2 DVSS 0.141794f
C1812 a_6164_n9984.n3 DVSS 0.27805f
C1813 a_6164_n9984.t13 DVSS 0.049102f
C1814 a_6164_n9984.t12 DVSS 0.049102f
C1815 a_6164_n9984.n4 DVSS 0.141794f
C1816 a_6164_n9984.n5 DVSS 0.27805f
C1817 a_6164_n9984.t7 DVSS 0.049102f
C1818 a_6164_n9984.t6 DVSS 0.049102f
C1819 a_6164_n9984.n6 DVSS 0.141794f
C1820 a_6164_n9984.n7 DVSS 0.27805f
C1821 a_6164_n9984.t14 DVSS 0.049102f
C1822 a_6164_n9984.t17 DVSS 0.049102f
C1823 a_6164_n9984.n8 DVSS 0.141794f
C1824 a_6164_n9984.n9 DVSS 0.278204f
C1825 a_6164_n9984.t8 DVSS 0.049102f
C1826 a_6164_n9984.t15 DVSS 0.049102f
C1827 a_6164_n9984.n10 DVSS 0.141794f
C1828 a_6164_n9984.n11 DVSS 0.370602f
C1829 a_6164_n9984.t9 DVSS 0.171712f
C1830 a_6164_n9984.n12 DVSS 0.519358f
C1831 a_6164_n9984.t27 DVSS 0.077863f
C1832 a_6164_n9984.n13 DVSS 1.07841f
C1833 a_6164_n9984.t20 DVSS 0.077863f
C1834 a_6164_n9984.n14 DVSS 0.761849f
C1835 a_6164_n9984.t25 DVSS 0.077863f
C1836 a_6164_n9984.n15 DVSS 0.761849f
C1837 a_6164_n9984.t1 DVSS 0.077863f
C1838 a_6164_n9984.n16 DVSS 0.761849f
C1839 a_6164_n9984.t3 DVSS 0.077863f
C1840 a_6164_n9984.n17 DVSS 0.761849f
C1841 a_6164_n9984.t2 DVSS 0.077863f
C1842 a_6164_n9984.n18 DVSS 0.761849f
C1843 a_6164_n9984.t18 DVSS 0.077863f
C1844 a_6164_n9984.n19 DVSS 0.761849f
C1845 a_6164_n9984.t22 DVSS 0.077863f
C1846 a_6164_n9984.n20 DVSS 0.761849f
C1847 a_6164_n9984.t19 DVSS 0.077863f
C1848 a_6164_n9984.n21 DVSS 0.761849f
C1849 a_6164_n9984.t24 DVSS 0.077863f
C1850 a_6164_n9984.n22 DVSS 0.761849f
C1851 a_6164_n9984.t29 DVSS 0.077863f
C1852 a_6164_n9984.n23 DVSS 0.761849f
C1853 a_6164_n9984.t28 DVSS 0.077863f
C1854 a_6164_n9984.n24 DVSS 0.761849f
C1855 a_6164_n9984.t21 DVSS 0.077863f
C1856 a_6164_n9984.n25 DVSS 0.761849f
C1857 a_6164_n9984.t23 DVSS 0.08f
C1858 a_6164_n9984.t26 DVSS 0.077863f
C1859 a_6164_n9984.n26 DVSS 1.42878f
C1860 a_6164_n9984.n27 DVSS 0.494727f
C1861 a_6164_n9984.t0 DVSS 0.344984f
C1862 D43v3.n0 DVSS 10.7802f
C1863 D43v3.n1 DVSS 10.7802f
C1864 D43v3.n2 DVSS 6.20209f
C1865 D43v3.n3 DVSS 6.6818f
C1866 D43v3.t0 DVSS 0.036168f
C1867 D43v3.t19 DVSS 0.821144f
C1868 D43v3.t21 DVSS 0.816878f
C1869 D43v3.t7 DVSS 0.816878f
C1870 D43v3.t9 DVSS 0.816878f
C1871 D43v3.t3 DVSS 0.816878f
C1872 D43v3.t23 DVSS 0.816878f
C1873 D43v3.t25 DVSS 0.816878f
C1874 D43v3.t11 DVSS 0.816878f
C1875 D43v3.t13 DVSS 0.816878f
C1876 D43v3.t5 DVSS 0.816878f
C1877 D43v3.t27 DVSS 0.816878f
C1878 D43v3.t29 DVSS 0.816878f
C1879 D43v3.t15 DVSS 0.816878f
C1880 D43v3.t17 DVSS 0.766841f
C1881 D43v3.t16 DVSS 0.766922f
C1882 D43v3.t18 DVSS 0.821144f
C1883 D43v3.t20 DVSS 0.816878f
C1884 D43v3.t6 DVSS 0.816878f
C1885 D43v3.t8 DVSS 0.816878f
C1886 D43v3.t2 DVSS 0.816878f
C1887 D43v3.t22 DVSS 0.816878f
C1888 D43v3.t24 DVSS 0.816878f
C1889 D43v3.t10 DVSS 0.816878f
C1890 D43v3.t12 DVSS 0.816878f
C1891 D43v3.t4 DVSS 0.816878f
C1892 D43v3.t26 DVSS 0.816878f
C1893 D43v3.t28 DVSS 0.816878f
C1894 D43v3.t14 DVSS 0.816878f
C1895 D43v3.n4 DVSS 2.63555f
C1896 D43v3.n5 DVSS 2.51841f
C1897 D43v3.n6 DVSS 0.030505f
C1898 D43v3.t1 DVSS 0.033965f
C1899 D43v3.n7 DVSS 0.029962f
C1900 x4.V2.t92 DVSS 0.156749f
C1901 x4.V2.t79 DVSS 0.039813f
C1902 x4.V2.t76 DVSS 0.039813f
C1903 x4.V2.n0 DVSS 0.131671f
C1904 x4.V2.t85 DVSS 0.039813f
C1905 x4.V2.t9 DVSS 0.039813f
C1906 x4.V2.n1 DVSS 0.123823f
C1907 x4.V2.n2 DVSS 0.408766f
C1908 x4.V2.t5 DVSS 0.039813f
C1909 x4.V2.t77 DVSS 0.039813f
C1910 x4.V2.n3 DVSS 0.123823f
C1911 x4.V2.n4 DVSS 0.233692f
C1912 x4.V2.t11 DVSS 0.039813f
C1913 x4.V2.t10 DVSS 0.039813f
C1914 x4.V2.n5 DVSS 0.123823f
C1915 x4.V2.n6 DVSS 0.233692f
C1916 x4.V2.t63 DVSS 0.039813f
C1917 x4.V2.t6 DVSS 0.039813f
C1918 x4.V2.n7 DVSS 0.123823f
C1919 x4.V2.n8 DVSS 0.23358f
C1920 x4.V2.t22 DVSS 0.039813f
C1921 x4.V2.t23 DVSS 0.039813f
C1922 x4.V2.n9 DVSS 0.123823f
C1923 x4.V2.n10 DVSS 0.23358f
C1924 x4.V2.t83 DVSS 0.039813f
C1925 x4.V2.t84 DVSS 0.039813f
C1926 x4.V2.n11 DVSS 0.123823f
C1927 x4.V2.n12 DVSS 0.276376f
C1928 x4.V2.t61 DVSS 0.039632f
C1929 x4.V2.t17 DVSS 0.039632f
C1930 x4.V2.n13 DVSS 0.123166f
C1931 x4.V2.n14 DVSS 0.275785f
C1932 x4.V2.t19 DVSS 0.039632f
C1933 x4.V2.t18 DVSS 0.039632f
C1934 x4.V2.n15 DVSS 0.123166f
C1935 x4.V2.n16 DVSS 0.23299f
C1936 x4.V2.t62 DVSS 0.039632f
C1937 x4.V2.t42 DVSS 0.039632f
C1938 x4.V2.n17 DVSS 0.123166f
C1939 x4.V2.n18 DVSS 0.23299f
C1940 x4.V2.t43 DVSS 0.039632f
C1941 x4.V2.t60 DVSS 0.039632f
C1942 x4.V2.n19 DVSS 0.123166f
C1943 x4.V2.n20 DVSS 0.275785f
C1944 x4.V2.t34 DVSS 0.042075f
C1945 x4.V2.t36 DVSS 0.042075f
C1946 x4.V2.n21 DVSS 0.131917f
C1947 x4.V2.n22 DVSS 0.285287f
C1948 x4.V2.t25 DVSS 0.042075f
C1949 x4.V2.t35 DVSS 0.042075f
C1950 x4.V2.n23 DVSS 0.131917f
C1951 x4.V2.n24 DVSS 0.285287f
C1952 x4.V2.t40 DVSS 0.044065f
C1953 x4.V2.t41 DVSS 0.044065f
C1954 x4.V2.n25 DVSS 0.141937f
C1955 x4.V2.n26 DVSS 0.332914f
C1956 x4.V2.t59 DVSS 0.196844f
C1957 x4.V2.n27 DVSS 0.371104f
C1958 x4.V2.n28 DVSS 0.243863f
C1959 x4.V2.t94 DVSS 1.63641f
C1960 x4.V2.n29 DVSS 0.291818f
C1961 x4.V2.t64 DVSS 0.064521f
C1962 x4.V2.n30 DVSS 0.648014f
C1963 x4.V2.t28 DVSS 0.051622f
C1964 x4.V2.n31 DVSS 0.449793f
C1965 x4.V2.t58 DVSS 0.051622f
C1966 x4.V2.n32 DVSS 0.315406f
C1967 x4.V2.t12 DVSS 0.051622f
C1968 x4.V2.n33 DVSS 0.449793f
C1969 x4.V2.t57 DVSS 0.051622f
C1970 x4.V2.n34 DVSS 0.315406f
C1971 x4.V2.t71 DVSS 0.051622f
C1972 x4.V2.n35 DVSS 0.449793f
C1973 x4.V2.t72 DVSS 0.051622f
C1974 x4.V2.n36 DVSS 0.315406f
C1975 x4.V2.t69 DVSS 0.051622f
C1976 x4.V2.n37 DVSS 0.449793f
C1977 x4.V2.n38 DVSS 0.315406f
C1978 x4.V2.t1 DVSS 0.051622f
C1979 x4.V2.n39 DVSS 0.449793f
C1980 x4.V2.t27 DVSS 0.051622f
C1981 x4.V2.n40 DVSS 0.315406f
C1982 x4.V2.t65 DVSS 0.051622f
C1983 x4.V2.n41 DVSS 0.449793f
C1984 x4.V2.t3 DVSS 0.051622f
C1985 x4.V2.n42 DVSS 0.315406f
C1986 x4.V2.t66 DVSS 0.051622f
C1987 x4.V2.n43 DVSS 0.449793f
C1988 x4.V2.t37 DVSS 0.051622f
C1989 x4.V2.n44 DVSS 0.315406f
C1990 x4.V2.t91 DVSS 0.051622f
C1991 x4.V2.n45 DVSS 0.449793f
C1992 x4.V2.t20 DVSS 0.051622f
C1993 x4.V2.n46 DVSS 0.315406f
C1994 x4.V2.t46 DVSS 0.051622f
C1995 x4.V2.n47 DVSS 0.449793f
C1996 x4.V2.t29 DVSS 0.051622f
C1997 x4.V2.n48 DVSS 0.315406f
C1998 x4.V2.t50 DVSS 0.051622f
C1999 x4.V2.n49 DVSS 0.449793f
C2000 x4.V2.t82 DVSS 0.051622f
C2001 x4.V2.n50 DVSS 0.315406f
C2002 x4.V2.t78 DVSS 0.051622f
C2003 x4.V2.n51 DVSS 0.449793f
C2004 x4.V2.t38 DVSS 0.051622f
C2005 x4.V2.n52 DVSS 0.315406f
C2006 x4.V2.t80 DVSS 0.051622f
C2007 x4.V2.n53 DVSS 0.449793f
C2008 x4.V2.t51 DVSS 0.051622f
C2009 x4.V2.n54 DVSS 0.315406f
C2010 x4.V2.t49 DVSS 0.051622f
C2011 x4.V2.n55 DVSS 0.449793f
C2012 x4.V2.t87 DVSS 0.051622f
C2013 x4.V2.n56 DVSS 0.315406f
C2014 x4.V2.t52 DVSS 0.051622f
C2015 x4.V2.n57 DVSS 0.449793f
C2016 x4.V2.t75 DVSS 0.051622f
C2017 x4.V2.t13 DVSS 0.051622f
C2018 x4.V2.n58 DVSS 0.449793f
C2019 x4.V2.t56 DVSS 0.272224f
C2020 x4.V2.t45 DVSS 0.186009f
C2021 x4.V2.n59 DVSS 0.169897f
C2022 x4.V2.t54 DVSS 0.186009f
C2023 x4.V2.n60 DVSS 0.160405f
C2024 x4.V2.t88 DVSS 0.186009f
C2025 x4.V2.n61 DVSS 0.160405f
C2026 x4.V2.t89 DVSS 0.051622f
C2027 x4.V2.n62 DVSS 0.457306f
C2028 x4.V2.n63 DVSS 0.187975f
C2029 x4.V2.n64 DVSS 0.528835f
C2030 x4.V2.n65 DVSS 0.315406f
C2031 x4.V2.n66 DVSS 0.449793f
C2032 x4.V2.t2 DVSS 0.051622f
C2033 x4.V2.n67 DVSS 0.449793f
C2034 x4.V2.t67 DVSS 0.051622f
C2035 x4.V2.n68 DVSS 0.449793f
C2036 x4.V2.n69 DVSS 0.315406f
C2037 x4.V2.n70 DVSS 0.315406f
C2038 x4.V2.n71 DVSS 0.315406f
C2039 x4.V2.n72 DVSS 0.449793f
C2040 x4.V2.t4 DVSS 0.051622f
C2041 x4.V2.n73 DVSS 0.449793f
C2042 x4.V2.t15 DVSS 0.051622f
C2043 x4.V2.n74 DVSS 0.449793f
C2044 x4.V2.n75 DVSS 0.315406f
C2045 x4.V2.n76 DVSS 0.315406f
C2046 x4.V2.n77 DVSS 0.315406f
C2047 x4.V2.n78 DVSS 0.449793f
C2048 x4.V2.t48 DVSS 0.051622f
C2049 x4.V2.n79 DVSS 0.449793f
C2050 x4.V2.t93 DVSS 0.051622f
C2051 x4.V2.n80 DVSS 0.449793f
C2052 x4.V2.n81 DVSS 0.315406f
C2053 x4.V2.n82 DVSS 0.315406f
C2054 x4.V2.n83 DVSS 0.315406f
C2055 x4.V2.n84 DVSS 0.449793f
C2056 x4.V2.t44 DVSS 0.051622f
C2057 x4.V2.n85 DVSS 0.449793f
C2058 x4.V2.t21 DVSS 0.051622f
C2059 x4.V2.n86 DVSS 0.449793f
C2060 x4.V2.n87 DVSS 0.315406f
C2061 x4.V2.n88 DVSS 0.315406f
C2062 x4.V2.n89 DVSS 0.315406f
C2063 x4.V2.n90 DVSS 0.449793f
C2064 x4.V2.t90 DVSS 0.051622f
C2065 x4.V2.n91 DVSS 0.449793f
C2066 x4.V2.t8 DVSS 0.051622f
C2067 x4.V2.n92 DVSS 0.449793f
C2068 x4.V2.n93 DVSS 0.315406f
C2069 x4.V2.n94 DVSS 0.315406f
C2070 x4.V2.n95 DVSS 0.315406f
C2071 x4.V2.n96 DVSS 0.449793f
C2072 x4.V2.t55 DVSS 0.051622f
C2073 x4.V2.n97 DVSS 0.449793f
C2074 x4.V2.t30 DVSS 0.051622f
C2075 x4.V2.n98 DVSS 0.449793f
C2076 x4.V2.n99 DVSS 0.315406f
C2077 x4.V2.n100 DVSS 0.315406f
C2078 x4.V2.n101 DVSS 0.315406f
C2079 x4.V2.n102 DVSS 0.449793f
C2080 x4.V2.t68 DVSS 0.051622f
C2081 x4.V2.n103 DVSS 0.449793f
C2082 x4.V2.t39 DVSS 0.051622f
C2083 x4.V2.n104 DVSS 0.449793f
C2084 x4.V2.n105 DVSS 0.315406f
C2085 x4.V2.n106 DVSS 0.315406f
C2086 x4.V2.n107 DVSS 0.315406f
C2087 x4.V2.n108 DVSS 0.449793f
C2088 x4.V2.t70 DVSS 0.051622f
C2089 x4.V2.n109 DVSS 0.449793f
C2090 x4.V2.t33 DVSS 0.051622f
C2091 x4.V2.n110 DVSS 0.449793f
C2092 x4.V2.n111 DVSS 0.315406f
C2093 x4.V2.n112 DVSS 0.315406f
C2094 x4.V2.n113 DVSS 0.315406f
C2095 x4.V2.n114 DVSS 0.449793f
C2096 x4.V2.t26 DVSS 0.051622f
C2097 x4.V2.n115 DVSS 0.449793f
C2098 x4.V2.t32 DVSS 0.051622f
C2099 x4.V2.n116 DVSS 0.449793f
C2100 x4.V2.n117 DVSS 0.315406f
C2101 x4.V2.n118 DVSS 0.315406f
C2102 x4.V2.n119 DVSS 0.315406f
C2103 x4.V2.n120 DVSS 0.449793f
C2104 x4.V2.t47 DVSS 0.051622f
C2105 x4.V2.n121 DVSS 0.449793f
C2106 x4.V2.t31 DVSS 0.051622f
C2107 x4.V2.n122 DVSS 0.449793f
C2108 x4.V2.n123 DVSS 0.315406f
C2109 x4.V2.n124 DVSS 0.315406f
C2110 x4.V2.n125 DVSS 0.315406f
C2111 x4.V2.t0 DVSS 0.186009f
C2112 x4.V2.n126 DVSS 0.315406f
C2113 x4.V2.t81 DVSS 0.051622f
C2114 x4.V2.n127 DVSS 0.449793f
C2115 x4.V2.t73 DVSS 0.051622f
C2116 x4.V2.n128 DVSS 0.449793f
C2117 x4.V2.n129 DVSS 0.315406f
C2118 x4.V2.n130 DVSS 0.315406f
C2119 x4.V2.n131 DVSS 0.315406f
C2120 x4.V2.n132 DVSS 0.449793f
C2121 x4.V2.t74 DVSS 0.051622f
C2122 x4.V2.n133 DVSS 0.449793f
C2123 x4.V2.t16 DVSS 0.051622f
C2124 x4.V2.n134 DVSS 0.449793f
C2125 x4.V2.n135 DVSS 0.315406f
C2126 x4.V2.n136 DVSS 0.315406f
C2127 x4.V2.n137 DVSS 0.315406f
C2128 x4.V2.n138 DVSS 0.449793f
C2129 x4.V2.t86 DVSS 0.051622f
C2130 x4.V2.n139 DVSS 0.449793f
C2131 x4.V2.t53 DVSS 0.051622f
C2132 x4.V2.n140 DVSS 0.449793f
C2133 x4.V2.n141 DVSS 0.315406f
C2134 x4.V2.n142 DVSS 0.315406f
C2135 x4.V2.n143 DVSS 0.315406f
C2136 x4.V2.n144 DVSS 0.449793f
C2137 x4.V2.t14 DVSS 0.051622f
C2138 x4.V2.n145 DVSS 0.449793f
C2139 x4.V2.t7 DVSS 0.051622f
C2140 x4.V2.t24 DVSS 0.051622f
C2141 x4.V2.n146 DVSS 0.449793f
C2142 x4.V2.n147 DVSS 0.449793f
C2143 x4.V2.n148 DVSS 0.471587f
C2144 x4.V2.n149 DVSS 1.76612f
C2145 x4.V2.n150 DVSS 1.27681f
C2146 x4.V2.n151 DVSS 2.40269f
C2147 x5.V2.t77 DVSS 0.037074f
C2148 x5.V2.t78 DVSS 0.037074f
C2149 x5.V2.n0 DVSS 0.122614f
C2150 x5.V2.t83 DVSS 0.037074f
C2151 x5.V2.t84 DVSS 0.037074f
C2152 x5.V2.n1 DVSS 0.115306f
C2153 x5.V2.n2 DVSS 0.380648f
C2154 x5.V2.t47 DVSS 0.037074f
C2155 x5.V2.t75 DVSS 0.037074f
C2156 x5.V2.n3 DVSS 0.115306f
C2157 x5.V2.n4 DVSS 0.217617f
C2158 x5.V2.t9 DVSS 0.037074f
C2159 x5.V2.t8 DVSS 0.037074f
C2160 x5.V2.n5 DVSS 0.115306f
C2161 x5.V2.n6 DVSS 0.217617f
C2162 x5.V2.t61 DVSS 0.037074f
C2163 x5.V2.t5 DVSS 0.037074f
C2164 x5.V2.n7 DVSS 0.115306f
C2165 x5.V2.n8 DVSS 0.217513f
C2166 x5.V2.t10 DVSS 0.037074f
C2167 x5.V2.t21 DVSS 0.037074f
C2168 x5.V2.n9 DVSS 0.115306f
C2169 x5.V2.n10 DVSS 0.217513f
C2170 x5.V2.t62 DVSS 0.037074f
C2171 x5.V2.t82 DVSS 0.037074f
C2172 x5.V2.n11 DVSS 0.115306f
C2173 x5.V2.n12 DVSS 0.257364f
C2174 x5.V2.t58 DVSS 0.036906f
C2175 x5.V2.t16 DVSS 0.036906f
C2176 x5.V2.n13 DVSS 0.114693f
C2177 x5.V2.n14 DVSS 0.256815f
C2178 x5.V2.t18 DVSS 0.036906f
C2179 x5.V2.t60 DVSS 0.036906f
C2180 x5.V2.n15 DVSS 0.114693f
C2181 x5.V2.n16 DVSS 0.216963f
C2182 x5.V2.t59 DVSS 0.036906f
C2183 x5.V2.t17 DVSS 0.036906f
C2184 x5.V2.n17 DVSS 0.114693f
C2185 x5.V2.n18 DVSS 0.216963f
C2186 x5.V2.t41 DVSS 0.036906f
C2187 x5.V2.t26 DVSS 0.036906f
C2188 x5.V2.n19 DVSS 0.114693f
C2189 x5.V2.n20 DVSS 0.206466f
C2190 x5.V2.t92 DVSS 0.145966f
C2191 x5.V2.n21 DVSS 0.227088f
C2192 x5.V2.t34 DVSS 0.183303f
C2193 x5.V2.n22 DVSS 0.345577f
C2194 x5.V2.t91 DVSS 0.041034f
C2195 x5.V2.t40 DVSS 0.041034f
C2196 x5.V2.n23 DVSS 0.132173f
C2197 x5.V2.n24 DVSS 0.310014f
C2198 x5.V2.t23 DVSS 0.039181f
C2199 x5.V2.t25 DVSS 0.039181f
C2200 x5.V2.n25 DVSS 0.122842f
C2201 x5.V2.n26 DVSS 0.265663f
C2202 x5.V2.t24 DVSS 0.039181f
C2203 x5.V2.t36 DVSS 0.039181f
C2204 x5.V2.n27 DVSS 0.122842f
C2205 x5.V2.n28 DVSS 0.220759f
C2206 x5.V2.n29 DVSS 2.33447f
C2207 x5.V2.t94 DVSS 1.52385f
C2208 x5.V2.n30 DVSS 0.183255f
C2209 x5.V2.n31 DVSS 0.29371f
C2210 x5.V2.t32 DVSS 0.047894f
C2211 x5.V2.n32 DVSS 0.41903f
C2212 x5.V2.n33 DVSS 0.29371f
C2213 x5.V2.t33 DVSS 0.047894f
C2214 x5.V2.n34 DVSS 0.41903f
C2215 x5.V2.n35 DVSS 0.29371f
C2216 x5.V2.t35 DVSS 0.047894f
C2217 x5.V2.n36 DVSS 0.41903f
C2218 x5.V2.n37 DVSS 0.29371f
C2219 x5.V2.t39 DVSS 0.047894f
C2220 x5.V2.n38 DVSS 0.41903f
C2221 x5.V2.n39 DVSS 0.29371f
C2222 x5.V2.t31 DVSS 0.047894f
C2223 x5.V2.n40 DVSS 0.41903f
C2224 x5.V2.n41 DVSS 0.29371f
C2225 x5.V2.t7 DVSS 0.047894f
C2226 x5.V2.n42 DVSS 0.41903f
C2227 x5.V2.n43 DVSS 0.29371f
C2228 x5.V2.t20 DVSS 0.047894f
C2229 x5.V2.n44 DVSS 0.41903f
C2230 x5.V2.n45 DVSS 0.29371f
C2231 x5.V2.t93 DVSS 0.047894f
C2232 x5.V2.n46 DVSS 0.41903f
C2233 x5.V2.n47 DVSS 0.29371f
C2234 x5.V2.t14 DVSS 0.047894f
C2235 x5.V2.n48 DVSS 0.41903f
C2236 x5.V2.n49 DVSS 0.29371f
C2237 x5.V2.t66 DVSS 0.047894f
C2238 x5.V2.n50 DVSS 0.41903f
C2239 x5.V2.n51 DVSS 0.29371f
C2240 x5.V2.t12 DVSS 0.047894f
C2241 x5.V2.n52 DVSS 0.41903f
C2242 x5.V2.t55 DVSS 0.101689f
C2243 x5.V2.t43 DVSS 0.047898f
C2244 x5.V2.n53 DVSS 0.435335f
C2245 x5.V2.t53 DVSS 0.047898f
C2246 x5.V2.n54 DVSS 0.274687f
C2247 x5.V2.t87 DVSS 0.047898f
C2248 x5.V2.n55 DVSS 0.274687f
C2249 x5.V2.t88 DVSS 0.047894f
C2250 x5.V2.n56 DVSS 0.426027f
C2251 x5.V2.n57 DVSS 0.175045f
C2252 x5.V2.n58 DVSS 0.492458f
C2253 x5.V2.t51 DVSS 0.047894f
C2254 x5.V2.n59 DVSS 0.41903f
C2255 x5.V2.t74 DVSS 0.047894f
C2256 x5.V2.n60 DVSS 0.41903f
C2257 x5.V2.t2 DVSS 0.047894f
C2258 x5.V2.n61 DVSS 0.41903f
C2259 x5.V2.n62 DVSS 0.29371f
C2260 x5.V2.n63 DVSS 0.29371f
C2261 x5.V2.n64 DVSS 0.29371f
C2262 x5.V2.t48 DVSS 0.047894f
C2263 x5.V2.n65 DVSS 0.41903f
C2264 x5.V2.t86 DVSS 0.047894f
C2265 x5.V2.n66 DVSS 0.41903f
C2266 x5.V2.t4 DVSS 0.047894f
C2267 x5.V2.n67 DVSS 0.41903f
C2268 x5.V2.n68 DVSS 0.29371f
C2269 x5.V2.n69 DVSS 0.29371f
C2270 x5.V2.n70 DVSS 0.29371f
C2271 x5.V2.t79 DVSS 0.047894f
C2272 x5.V2.n71 DVSS 0.41903f
C2273 x5.V2.t50 DVSS 0.047894f
C2274 x5.V2.n72 DVSS 0.41903f
C2275 x5.V2.t46 DVSS 0.047894f
C2276 x5.V2.n73 DVSS 0.41903f
C2277 x5.V2.n74 DVSS 0.29371f
C2278 x5.V2.n75 DVSS 0.29371f
C2279 x5.V2.n76 DVSS 0.29371f
C2280 x5.V2.t76 DVSS 0.047894f
C2281 x5.V2.n77 DVSS 0.41903f
C2282 x5.V2.t38 DVSS 0.047894f
C2283 x5.V2.n78 DVSS 0.41903f
C2284 x5.V2.t42 DVSS 0.047894f
C2285 x5.V2.n79 DVSS 0.41903f
C2286 x5.V2.n80 DVSS 0.29371f
C2287 x5.V2.n81 DVSS 0.29371f
C2288 x5.V2.n82 DVSS 0.29371f
C2289 x5.V2.t49 DVSS 0.047894f
C2290 x5.V2.n83 DVSS 0.41903f
C2291 x5.V2.t81 DVSS 0.047894f
C2292 x5.V2.n84 DVSS 0.41903f
C2293 x5.V2.t89 DVSS 0.047894f
C2294 x5.V2.n85 DVSS 0.41903f
C2295 x5.V2.n86 DVSS 0.29371f
C2296 x5.V2.n87 DVSS 0.29371f
C2297 x5.V2.n88 DVSS 0.29371f
C2298 x5.V2.t44 DVSS 0.047894f
C2299 x5.V2.n89 DVSS 0.41903f
C2300 x5.V2.t30 DVSS 0.047894f
C2301 x5.V2.n90 DVSS 0.41903f
C2302 x5.V2.t54 DVSS 0.047894f
C2303 x5.V2.n91 DVSS 0.41903f
C2304 x5.V2.n92 DVSS 0.29371f
C2305 x5.V2.n93 DVSS 0.29371f
C2306 x5.V2.n94 DVSS 0.29371f
C2307 x5.V2.t90 DVSS 0.047894f
C2308 x5.V2.n95 DVSS 0.41903f
C2309 x5.V2.t19 DVSS 0.047894f
C2310 x5.V2.n96 DVSS 0.41903f
C2311 x5.V2.t67 DVSS 0.047894f
C2312 x5.V2.n97 DVSS 0.41903f
C2313 x5.V2.n98 DVSS 0.29371f
C2314 x5.V2.n99 DVSS 0.29371f
C2315 x5.V2.n100 DVSS 0.29371f
C2316 x5.V2.t65 DVSS 0.047894f
C2317 x5.V2.n101 DVSS 0.41903f
C2318 x5.V2.t37 DVSS 0.047894f
C2319 x5.V2.n102 DVSS 0.41903f
C2320 x5.V2.t69 DVSS 0.047894f
C2321 x5.V2.n103 DVSS 0.41903f
C2322 x5.V2.n104 DVSS 0.29371f
C2323 x5.V2.n105 DVSS 0.29371f
C2324 x5.V2.n106 DVSS 0.29371f
C2325 x5.V2.t64 DVSS 0.047894f
C2326 x5.V2.n107 DVSS 0.41903f
C2327 x5.V2.t3 DVSS 0.047894f
C2328 x5.V2.n108 DVSS 0.41903f
C2329 x5.V2.t27 DVSS 0.047894f
C2330 x5.V2.n109 DVSS 0.41903f
C2331 x5.V2.n110 DVSS 0.29371f
C2332 x5.V2.n111 DVSS 0.29371f
C2333 x5.V2.n112 DVSS 0.29371f
C2334 x5.V2.t1 DVSS 0.047894f
C2335 x5.V2.n113 DVSS 0.41903f
C2336 x5.V2.t28 DVSS 0.047894f
C2337 x5.V2.n114 DVSS 0.41903f
C2338 x5.V2.t45 DVSS 0.047894f
C2339 x5.V2.n115 DVSS 0.41903f
C2340 x5.V2.n116 DVSS 0.29371f
C2341 x5.V2.n117 DVSS 0.29371f
C2342 x5.V2.n118 DVSS 0.29371f
C2343 x5.V2.t68 DVSS 0.047894f
C2344 x5.V2.n119 DVSS 0.41903f
C2345 x5.V2.t0 DVSS 0.047898f
C2346 x5.V2.n120 DVSS 0.419026f
C2347 x5.V2.t71 DVSS 0.047894f
C2348 x5.V2.n121 DVSS 0.41903f
C2349 x5.V2.n122 DVSS 0.29371f
C2350 x5.V2.t56 DVSS 0.047894f
C2351 x5.V2.n123 DVSS 0.41903f
C2352 x5.V2.n124 DVSS 0.29371f
C2353 x5.V2.t57 DVSS 0.047894f
C2354 x5.V2.n125 DVSS 0.41903f
C2355 x5.V2.n126 DVSS 0.564037f
C2356 x5.V2.t63 DVSS 0.059963f
C2357 x5.V2.n127 DVSS 0.603559f
C2358 x5.V2.t22 DVSS 0.047894f
C2359 x5.V2.n128 DVSS 0.41903f
C2360 x5.V2.t6 DVSS 0.047894f
C2361 x5.V2.n129 DVSS 0.41903f
C2362 x5.V2.t13 DVSS 0.047894f
C2363 x5.V2.n130 DVSS 0.41903f
C2364 x5.V2.n131 DVSS 0.29371f
C2365 x5.V2.n132 DVSS 0.29371f
C2366 x5.V2.n133 DVSS 0.29371f
C2367 x5.V2.t29 DVSS 0.047894f
C2368 x5.V2.n134 DVSS 0.41903f
C2369 x5.V2.t52 DVSS 0.047894f
C2370 x5.V2.n135 DVSS 0.41903f
C2371 x5.V2.t85 DVSS 0.047894f
C2372 x5.V2.n136 DVSS 0.41903f
C2373 x5.V2.n137 DVSS 0.29371f
C2374 x5.V2.n138 DVSS 0.29371f
C2375 x5.V2.n139 DVSS 0.29371f
C2376 x5.V2.t11 DVSS 0.047894f
C2377 x5.V2.n140 DVSS 0.41903f
C2378 x5.V2.t15 DVSS 0.047894f
C2379 x5.V2.n141 DVSS 0.41903f
C2380 x5.V2.t73 DVSS 0.047894f
C2381 x5.V2.n142 DVSS 0.41903f
C2382 x5.V2.n143 DVSS 0.29371f
C2383 x5.V2.n144 DVSS 0.29371f
C2384 x5.V2.n145 DVSS 0.29371f
C2385 x5.V2.t70 DVSS 0.047894f
C2386 x5.V2.n146 DVSS 0.41903f
C2387 x5.V2.t72 DVSS 0.047894f
C2388 x5.V2.n147 DVSS 0.41903f
C2389 x5.V2.t80 DVSS 0.047894f
C2390 x5.V2.n148 DVSS 0.41903f
C2391 x5.V2.n149 DVSS 0.25731f
C2392 x5.V2.n150 DVSS 1.96593f
C2393 x5.V2.n151 DVSS 1.92469f
C2394 x5.V2.n152 DVSS 3.89658f
C2395 x3.R1.t74 DVSS 0.034323f
C2396 x3.R1.t72 DVSS 0.034323f
C2397 x3.R1.n0 DVSS 0.113516f
C2398 x3.R1.t78 DVSS 0.034323f
C2399 x3.R1.t79 DVSS 0.034323f
C2400 x3.R1.n1 DVSS 0.10675f
C2401 x3.R1.n2 DVSS 0.352403f
C2402 x3.R1.t67 DVSS 0.034323f
C2403 x3.R1.t71 DVSS 0.034323f
C2404 x3.R1.n3 DVSS 0.10675f
C2405 x3.R1.n4 DVSS 0.20147f
C2406 x3.R1.t70 DVSS 0.034323f
C2407 x3.R1.t77 DVSS 0.034323f
C2408 x3.R1.n5 DVSS 0.10675f
C2409 x3.R1.n6 DVSS 0.20147f
C2410 x3.R1.t76 DVSS 0.034323f
C2411 x3.R1.t66 DVSS 0.034323f
C2412 x3.R1.n7 DVSS 0.10675f
C2413 x3.R1.n8 DVSS 0.201373f
C2414 x3.R1.t69 DVSS 0.034323f
C2415 x3.R1.t68 DVSS 0.034323f
C2416 x3.R1.n9 DVSS 0.10675f
C2417 x3.R1.n10 DVSS 0.201373f
C2418 x3.R1.t75 DVSS 0.034323f
C2419 x3.R1.t73 DVSS 0.034323f
C2420 x3.R1.n11 DVSS 0.10675f
C2421 x3.R1.n12 DVSS 0.189509f
C2422 x3.R1.t92 DVSS 0.135135f
C2423 x3.R1.n13 DVSS 0.210238f
C2424 x3.R1.t26 DVSS 0.169702f
C2425 x3.R1.n14 DVSS 0.319935f
C2426 x3.R1.t55 DVSS 0.037989f
C2427 x3.R1.t56 DVSS 0.037989f
C2428 x3.R1.n15 DVSS 0.122366f
C2429 x3.R1.n16 DVSS 0.28701f
C2430 x3.R1.t16 DVSS 0.036273f
C2431 x3.R1.t15 DVSS 0.036273f
C2432 x3.R1.n17 DVSS 0.113727f
C2433 x3.R1.n18 DVSS 0.24595f
C2434 x3.R1.t18 DVSS 0.036273f
C2435 x3.R1.t8 DVSS 0.036273f
C2436 x3.R1.n19 DVSS 0.113727f
C2437 x3.R1.n20 DVSS 0.24595f
C2438 x3.R1.t59 DVSS 0.034167f
C2439 x3.R1.t62 DVSS 0.034167f
C2440 x3.R1.n21 DVSS 0.106183f
C2441 x3.R1.n22 DVSS 0.237759f
C2442 x3.R1.t64 DVSS 0.034167f
C2443 x3.R1.t58 DVSS 0.034167f
C2444 x3.R1.n23 DVSS 0.106183f
C2445 x3.R1.n24 DVSS 0.200864f
C2446 x3.R1.t65 DVSS 0.034167f
C2447 x3.R1.t42 DVSS 0.034167f
C2448 x3.R1.n25 DVSS 0.106183f
C2449 x3.R1.n26 DVSS 0.200864f
C2450 x3.R1.t63 DVSS 0.034167f
C2451 x3.R1.t60 DVSS 0.034167f
C2452 x3.R1.n27 DVSS 0.106183f
C2453 x3.R1.n28 DVSS 0.196463f
C2454 x3.R1.n29 DVSS 1.11035f
C2455 x3.R1.t94 DVSS 1.41114f
C2456 x3.R1.n30 DVSS 0.247514f
C2457 x3.R1.n31 DVSS 0.271917f
C2458 x3.R1.t90 DVSS 0.04434f
C2459 x3.R1.n32 DVSS 0.387938f
C2460 x3.R1.n33 DVSS 0.271917f
C2461 x3.R1.t37 DVSS 0.04434f
C2462 x3.R1.n34 DVSS 0.387938f
C2463 x3.R1.t0 DVSS 0.044344f
C2464 x3.R1.t24 DVSS 0.094144f
C2465 x3.R1.t36 DVSS 0.044344f
C2466 x3.R1.n35 DVSS 0.403033f
C2467 x3.R1.t82 DVSS 0.044344f
C2468 x3.R1.n36 DVSS 0.254305f
C2469 x3.R1.t35 DVSS 0.044344f
C2470 x3.R1.n37 DVSS 0.254305f
C2471 x3.R1.t31 DVSS 0.04434f
C2472 x3.R1.n38 DVSS 0.394415f
C2473 x3.R1.n39 DVSS 0.162056f
C2474 x3.R1.t29 DVSS 0.04434f
C2475 x3.R1.n40 DVSS 0.387938f
C2476 x3.R1.t14 DVSS 0.04434f
C2477 x3.R1.n41 DVSS 0.387938f
C2478 x3.R1.n42 DVSS 0.455917f
C2479 x3.R1.n43 DVSS 0.271917f
C2480 x3.R1.n44 DVSS 0.271917f
C2481 x3.R1.n45 DVSS 0.387934f
C2482 x3.R1.t46 DVSS 0.04434f
C2483 x3.R1.n46 DVSS 0.387938f
C2484 x3.R1.t57 DVSS 0.04434f
C2485 x3.R1.n47 DVSS 0.387938f
C2486 x3.R1.n48 DVSS 0.271917f
C2487 x3.R1.n49 DVSS 0.271917f
C2488 x3.R1.n50 DVSS 0.271917f
C2489 x3.R1.t83 DVSS 0.04434f
C2490 x3.R1.n51 DVSS 0.387938f
C2491 x3.R1.t11 DVSS 0.04434f
C2492 x3.R1.n52 DVSS 0.387938f
C2493 x3.R1.t2 DVSS 0.04434f
C2494 x3.R1.n53 DVSS 0.387938f
C2495 x3.R1.n54 DVSS 0.271917f
C2496 x3.R1.t28 DVSS 0.04434f
C2497 x3.R1.n55 DVSS 0.387938f
C2498 x3.R1.n56 DVSS 0.271917f
C2499 x3.R1.t85 DVSS 0.04434f
C2500 x3.R1.n57 DVSS 0.387938f
C2501 x3.R1.n58 DVSS 0.271917f
C2502 x3.R1.t41 DVSS 0.04434f
C2503 x3.R1.n59 DVSS 0.387938f
C2504 x3.R1.n60 DVSS 0.271917f
C2505 x3.R1.t5 DVSS 0.04434f
C2506 x3.R1.n61 DVSS 0.387938f
C2507 x3.R1.n62 DVSS 0.271917f
C2508 x3.R1.t81 DVSS 0.04434f
C2509 x3.R1.n63 DVSS 0.387938f
C2510 x3.R1.n64 DVSS 0.271917f
C2511 x3.R1.t89 DVSS 0.04434f
C2512 x3.R1.n65 DVSS 0.387938f
C2513 x3.R1.n66 DVSS 0.271917f
C2514 x3.R1.t23 DVSS 0.04434f
C2515 x3.R1.n67 DVSS 0.387938f
C2516 x3.R1.n68 DVSS 0.271917f
C2517 x3.R1.t87 DVSS 0.04434f
C2518 x3.R1.n69 DVSS 0.387938f
C2519 x3.R1.n70 DVSS 0.271917f
C2520 x3.R1.t32 DVSS 0.04434f
C2521 x3.R1.n71 DVSS 0.387938f
C2522 x3.R1.n72 DVSS 0.271917f
C2523 x3.R1.t51 DVSS 0.04434f
C2524 x3.R1.n73 DVSS 0.387938f
C2525 x3.R1.n74 DVSS 0.271917f
C2526 x3.R1.t44 DVSS 0.04434f
C2527 x3.R1.n75 DVSS 0.387938f
C2528 x3.R1.t53 DVSS 0.055514f
C2529 x3.R1.t48 DVSS 0.04434f
C2530 x3.R1.n76 DVSS 0.387938f
C2531 x3.R1.n77 DVSS 0.558774f
C2532 x3.R1.n78 DVSS 0.522185f
C2533 x3.R1.n79 DVSS 0.271917f
C2534 x3.R1.t93 DVSS 0.04434f
C2535 x3.R1.n80 DVSS 0.387938f
C2536 x3.R1.t9 DVSS 0.04434f
C2537 x3.R1.n81 DVSS 0.387938f
C2538 x3.R1.t20 DVSS 0.04434f
C2539 x3.R1.n82 DVSS 0.387938f
C2540 x3.R1.n83 DVSS 0.271917f
C2541 x3.R1.n84 DVSS 0.271917f
C2542 x3.R1.n85 DVSS 0.271917f
C2543 x3.R1.t38 DVSS 0.04434f
C2544 x3.R1.n86 DVSS 0.387938f
C2545 x3.R1.t22 DVSS 0.04434f
C2546 x3.R1.n87 DVSS 0.387938f
C2547 x3.R1.t27 DVSS 0.04434f
C2548 x3.R1.n88 DVSS 0.387938f
C2549 x3.R1.n89 DVSS 0.271917f
C2550 x3.R1.n90 DVSS 0.271917f
C2551 x3.R1.n91 DVSS 0.271917f
C2552 x3.R1.t4 DVSS 0.04434f
C2553 x3.R1.n92 DVSS 0.387938f
C2554 x3.R1.t17 DVSS 0.04434f
C2555 x3.R1.n93 DVSS 0.387938f
C2556 x3.R1.t84 DVSS 0.04434f
C2557 x3.R1.n94 DVSS 0.387938f
C2558 x3.R1.n95 DVSS 0.271917f
C2559 x3.R1.n96 DVSS 0.271917f
C2560 x3.R1.n97 DVSS 0.271917f
C2561 x3.R1.t19 DVSS 0.04434f
C2562 x3.R1.n98 DVSS 0.387938f
C2563 x3.R1.t33 DVSS 0.04434f
C2564 x3.R1.n99 DVSS 0.387938f
C2565 x3.R1.t54 DVSS 0.04434f
C2566 x3.R1.n100 DVSS 0.387938f
C2567 x3.R1.n101 DVSS 0.271917f
C2568 x3.R1.n102 DVSS 0.271917f
C2569 x3.R1.n103 DVSS 0.271917f
C2570 x3.R1.t1 DVSS 0.04434f
C2571 x3.R1.n104 DVSS 0.387938f
C2572 x3.R1.t91 DVSS 0.04434f
C2573 x3.R1.n105 DVSS 0.387938f
C2574 x3.R1.t40 DVSS 0.04434f
C2575 x3.R1.n106 DVSS 0.387938f
C2576 x3.R1.n107 DVSS 0.271917f
C2577 x3.R1.n108 DVSS 0.271917f
C2578 x3.R1.n109 DVSS 0.271917f
C2579 x3.R1.t47 DVSS 0.04434f
C2580 x3.R1.n110 DVSS 0.387938f
C2581 x3.R1.t80 DVSS 0.04434f
C2582 x3.R1.n111 DVSS 0.387938f
C2583 x3.R1.t6 DVSS 0.04434f
C2584 x3.R1.n112 DVSS 0.387938f
C2585 x3.R1.n113 DVSS 0.271917f
C2586 x3.R1.n114 DVSS 0.271917f
C2587 x3.R1.n115 DVSS 0.271917f
C2588 x3.R1.t7 DVSS 0.04434f
C2589 x3.R1.n116 DVSS 0.387938f
C2590 x3.R1.t39 DVSS 0.04434f
C2591 x3.R1.n117 DVSS 0.387938f
C2592 x3.R1.t88 DVSS 0.04434f
C2593 x3.R1.n118 DVSS 0.387938f
C2594 x3.R1.n119 DVSS 0.271917f
C2595 x3.R1.n120 DVSS 0.271917f
C2596 x3.R1.n121 DVSS 0.271917f
C2597 x3.R1.t45 DVSS 0.04434f
C2598 x3.R1.n122 DVSS 0.387938f
C2599 x3.R1.t25 DVSS 0.04434f
C2600 x3.R1.n123 DVSS 0.387938f
C2601 x3.R1.t12 DVSS 0.04434f
C2602 x3.R1.n124 DVSS 0.387938f
C2603 x3.R1.n125 DVSS 0.271917f
C2604 x3.R1.n126 DVSS 0.271917f
C2605 x3.R1.n127 DVSS 0.271917f
C2606 x3.R1.t86 DVSS 0.04434f
C2607 x3.R1.n128 DVSS 0.387938f
C2608 x3.R1.t43 DVSS 0.04434f
C2609 x3.R1.n129 DVSS 0.387938f
C2610 x3.R1.t21 DVSS 0.04434f
C2611 x3.R1.n130 DVSS 0.387938f
C2612 x3.R1.n131 DVSS 0.271917f
C2613 x3.R1.n132 DVSS 0.271917f
C2614 x3.R1.n133 DVSS 0.271917f
C2615 x3.R1.t52 DVSS 0.04434f
C2616 x3.R1.n134 DVSS 0.387938f
C2617 x3.R1.t3 DVSS 0.04434f
C2618 x3.R1.n135 DVSS 0.387938f
C2619 x3.R1.t50 DVSS 0.04434f
C2620 x3.R1.n136 DVSS 0.387938f
C2621 x3.R1.n137 DVSS 0.271917f
C2622 x3.R1.n138 DVSS 0.271917f
C2623 x3.R1.n139 DVSS 0.271917f
C2624 x3.R1.t34 DVSS 0.04434f
C2625 x3.R1.n140 DVSS 0.387938f
C2626 x3.R1.t61 DVSS 0.04434f
C2627 x3.R1.n141 DVSS 0.387938f
C2628 x3.R1.t10 DVSS 0.04434f
C2629 x3.R1.n142 DVSS 0.387938f
C2630 x3.R1.n143 DVSS 0.271917f
C2631 x3.R1.n144 DVSS 0.271917f
C2632 x3.R1.n145 DVSS 0.271917f
C2633 x3.R1.t30 DVSS 0.04434f
C2634 x3.R1.n146 DVSS 0.387938f
C2635 x3.R1.t49 DVSS 0.04434f
C2636 x3.R1.n147 DVSS 0.387938f
C2637 x3.R1.t13 DVSS 0.04434f
C2638 x3.R1.n148 DVSS 0.387938f
C2639 x3.R1.n149 DVSS 0.160361f
C2640 x3.R1.n150 DVSS 2.68934f
C2641 x3.R1.n151 DVSS 1.86014f
C2642 x3.R1.n152 DVSS 2.02828f
C2643 a_16261_n4916.t18 DVSS 0.213748f
C2644 a_16261_n4916.t25 DVSS 0.048284f
C2645 a_16261_n4916.t20 DVSS 0.048284f
C2646 a_16261_n4916.n0 DVSS 0.139431f
C2647 a_16261_n4916.n1 DVSS 0.50097f
C2648 a_16261_n4916.t23 DVSS 0.048284f
C2649 a_16261_n4916.t14 DVSS 0.048284f
C2650 a_16261_n4916.n2 DVSS 0.139431f
C2651 a_16261_n4916.n3 DVSS 0.273415f
C2652 a_16261_n4916.t22 DVSS 0.048284f
C2653 a_16261_n4916.t21 DVSS 0.048284f
C2654 a_16261_n4916.n4 DVSS 0.139431f
C2655 a_16261_n4916.n5 DVSS 0.273415f
C2656 a_16261_n4916.t16 DVSS 0.048284f
C2657 a_16261_n4916.t15 DVSS 0.048284f
C2658 a_16261_n4916.n6 DVSS 0.139431f
C2659 a_16261_n4916.n7 DVSS 0.273415f
C2660 a_16261_n4916.t27 DVSS 0.048284f
C2661 a_16261_n4916.t24 DVSS 0.048284f
C2662 a_16261_n4916.n8 DVSS 0.139431f
C2663 a_16261_n4916.n9 DVSS 0.273567f
C2664 a_16261_n4916.t17 DVSS 0.048284f
C2665 a_16261_n4916.t26 DVSS 0.048284f
C2666 a_16261_n4916.n10 DVSS 0.139431f
C2667 a_16261_n4916.n11 DVSS 0.364425f
C2668 a_16261_n4916.t19 DVSS 0.16885f
C2669 a_16261_n4916.n12 DVSS 0.510702f
C2670 a_16261_n4916.t28 DVSS 0.076565f
C2671 a_16261_n4916.n13 DVSS 1.06044f
C2672 a_16261_n4916.t6 DVSS 0.076565f
C2673 a_16261_n4916.n14 DVSS 0.749151f
C2674 a_16261_n4916.t7 DVSS 0.076565f
C2675 a_16261_n4916.n15 DVSS 0.749151f
C2676 a_16261_n4916.t29 DVSS 0.076565f
C2677 a_16261_n4916.n16 DVSS 0.749151f
C2678 a_16261_n4916.t4 DVSS 0.076565f
C2679 a_16261_n4916.n17 DVSS 0.749151f
C2680 a_16261_n4916.t8 DVSS 0.076565f
C2681 a_16261_n4916.n18 DVSS 0.749151f
C2682 a_16261_n4916.t13 DVSS 0.076565f
C2683 a_16261_n4916.n19 DVSS 0.749151f
C2684 a_16261_n4916.t3 DVSS 0.076565f
C2685 a_16261_n4916.n20 DVSS 0.749151f
C2686 a_16261_n4916.t9 DVSS 0.076565f
C2687 a_16261_n4916.n21 DVSS 0.749151f
C2688 a_16261_n4916.t10 DVSS 0.076565f
C2689 a_16261_n4916.n22 DVSS 0.749151f
C2690 a_16261_n4916.t11 DVSS 0.076565f
C2691 a_16261_n4916.n23 DVSS 0.749151f
C2692 a_16261_n4916.t2 DVSS 0.076565f
C2693 a_16261_n4916.n24 DVSS 0.749151f
C2694 a_16261_n4916.t12 DVSS 0.076565f
C2695 a_16261_n4916.n25 DVSS 0.749151f
C2696 a_16261_n4916.t5 DVSS 0.078667f
C2697 a_16261_n4916.t1 DVSS 0.076565f
C2698 a_16261_n4916.n26 DVSS 1.40496f
C2699 a_16261_n4916.n27 DVSS 0.486482f
C2700 a_16261_n4916.t0 DVSS 0.339234f
C2701 DVDD.n0 DVSS 0.071431f
C2702 DVDD.n1 DVSS 0.206741f
C2703 DVDD.t42 DVSS 0.270864f
C2704 DVDD.t24 DVSS 0.106135f
C2705 DVDD.n2 DVSS 0.095079f
C2706 DVDD.n4 DVSS 0.077524f
C2707 DVDD.n5 DVSS 0.118727f
C2708 DVDD.t43 DVSS 0.011257f
C2709 DVDD.t25 DVSS 0.011257f
C2710 DVDD.n6 DVSS 0.024688f
C2711 DVDD.n7 DVSS 0.320091f
C2712 DVDD.n8 DVSS 0.051683f
C2713 DVDD.n9 DVSS 0.027444f
C2714 DVDD.n10 DVSS 0.014242f
C2715 DVDD.t29 DVSS 0.011257f
C2716 DVDD.t37 DVSS 0.011257f
C2717 DVDD.n11 DVSS 0.024688f
C2718 DVDD.n12 DVSS 0.071431f
C2719 DVDD.n13 DVSS 0.206741f
C2720 DVDD.t28 DVSS 0.270864f
C2721 DVDD.t36 DVSS 0.106135f
C2722 DVDD.n14 DVSS 0.095079f
C2723 DVDD.n16 DVSS 0.077524f
C2724 DVDD.n17 DVSS 0.118727f
C2725 DVDD.t9 DVSS 0.011257f
C2726 DVDD.t1 DVSS 0.011257f
C2727 DVDD.n18 DVSS 0.024688f
C2728 DVDD.n19 DVSS 0.071431f
C2729 DVDD.n20 DVSS 0.206741f
C2730 DVDD.t8 DVSS 0.270864f
C2731 DVDD.t0 DVSS 0.106135f
C2732 DVDD.n21 DVSS 0.095079f
C2733 DVDD.n23 DVSS 0.077524f
C2734 DVDD.n24 DVSS 0.118727f
C2735 DVDD.t11 DVSS 0.011257f
C2736 DVDD.t7 DVSS 0.011257f
C2737 DVDD.n25 DVSS 0.024688f
C2738 DVDD.n26 DVSS 0.071431f
C2739 DVDD.n27 DVSS 0.206741f
C2740 DVDD.t10 DVSS 0.270864f
C2741 DVDD.t6 DVSS 0.106135f
C2742 DVDD.n28 DVSS 0.095079f
C2743 DVDD.n30 DVSS 0.077524f
C2744 DVDD.n31 DVSS 0.118727f
C2745 DVDD.t17 DVSS 0.011257f
C2746 DVDD.t13 DVSS 0.011257f
C2747 DVDD.n32 DVSS 0.024688f
C2748 DVDD.n33 DVSS 0.071431f
C2749 DVDD.n34 DVSS 0.206741f
C2750 DVDD.t16 DVSS 0.270864f
C2751 DVDD.t12 DVSS 0.106135f
C2752 DVDD.n35 DVSS 0.095079f
C2753 DVDD.n37 DVSS 0.077524f
C2754 DVDD.n38 DVSS 0.118727f
C2755 DVDD.t21 DVSS 0.011257f
C2756 DVDD.t35 DVSS 0.011257f
C2757 DVDD.n39 DVSS 0.024688f
C2758 DVDD.n40 DVSS 0.071431f
C2759 DVDD.n41 DVSS 0.206741f
C2760 DVDD.t20 DVSS 0.270864f
C2761 DVDD.t34 DVSS 0.106135f
C2762 DVDD.n42 DVSS 0.095079f
C2763 DVDD.n44 DVSS 0.077524f
C2764 DVDD.n45 DVSS 0.118727f
C2765 DVDD.t5 DVSS 0.011257f
C2766 DVDD.t41 DVSS 0.011257f
C2767 DVDD.n46 DVSS 0.024688f
C2768 DVDD.n47 DVSS 0.071431f
C2769 DVDD.n48 DVSS 0.206741f
C2770 DVDD.t4 DVSS 0.270864f
C2771 DVDD.t40 DVSS 0.106135f
C2772 DVDD.n49 DVSS 0.095079f
C2773 DVDD.n51 DVSS 0.077524f
C2774 DVDD.n52 DVSS 0.118727f
C2775 DVDD.t27 DVSS 0.011257f
C2776 DVDD.t19 DVSS 0.011257f
C2777 DVDD.n53 DVSS 0.024688f
C2778 DVDD.n54 DVSS 0.071431f
C2779 DVDD.n55 DVSS 0.206741f
C2780 DVDD.t26 DVSS 0.270864f
C2781 DVDD.t18 DVSS 0.106135f
C2782 DVDD.n56 DVSS 0.095079f
C2783 DVDD.n58 DVSS 0.077524f
C2784 DVDD.n59 DVSS 0.118727f
C2785 DVDD.t15 DVSS 0.011257f
C2786 DVDD.t39 DVSS 0.011257f
C2787 DVDD.n60 DVSS 0.024688f
C2788 DVDD.n61 DVSS 0.071431f
C2789 DVDD.n62 DVSS 0.206741f
C2790 DVDD.t14 DVSS 0.270864f
C2791 DVDD.t38 DVSS 0.106135f
C2792 DVDD.n63 DVSS 0.095079f
C2793 DVDD.n65 DVSS 0.077524f
C2794 DVDD.n66 DVSS 0.118727f
C2795 DVDD.t3 DVSS 0.011257f
C2796 DVDD.t23 DVSS 0.011257f
C2797 DVDD.n67 DVSS 0.024688f
C2798 DVDD.n68 DVSS 0.071431f
C2799 DVDD.n69 DVSS 0.206741f
C2800 DVDD.t2 DVSS 0.270864f
C2801 DVDD.t22 DVSS 0.106135f
C2802 DVDD.n70 DVSS 0.095079f
C2803 DVDD.n72 DVSS 0.077524f
C2804 DVDD.n73 DVSS 0.118727f
C2805 DVDD.t33 DVSS 0.011257f
C2806 DVDD.t31 DVSS 0.011257f
C2807 DVDD.n74 DVSS 0.024688f
C2808 DVDD.n75 DVSS 0.071431f
C2809 DVDD.n76 DVSS 0.206741f
C2810 DVDD.t32 DVSS 0.270864f
C2811 DVDD.t30 DVSS 0.106135f
C2812 DVDD.n77 DVSS 0.095079f
C2813 DVDD.n79 DVSS 0.077524f
C2814 DVDD.n80 DVSS 0.118727f
C2815 DVDD.n81 DVSS 0.014242f
C2816 DVDD.n82 DVSS 0.027444f
C2817 DVDD.n83 DVSS 0.051683f
C2818 DVDD.n84 DVSS 0.153995f
C2819 DVDD.n85 DVSS 0.014242f
C2820 DVDD.n86 DVSS 0.027444f
C2821 DVDD.n87 DVSS 0.051683f
C2822 DVDD.n88 DVSS 0.153995f
C2823 DVDD.n89 DVSS 0.014242f
C2824 DVDD.n90 DVSS 0.027444f
C2825 DVDD.n91 DVSS 0.051683f
C2826 DVDD.n92 DVSS 0.153995f
C2827 DVDD.n93 DVSS 0.014242f
C2828 DVDD.n94 DVSS 0.027444f
C2829 DVDD.n95 DVSS 0.051683f
C2830 DVDD.n96 DVSS 0.153995f
C2831 DVDD.n97 DVSS 0.014242f
C2832 DVDD.n98 DVSS 0.027444f
C2833 DVDD.n99 DVSS 0.051683f
C2834 DVDD.n100 DVSS 0.153995f
C2835 DVDD.n101 DVSS 0.014242f
C2836 DVDD.n102 DVSS 0.027444f
C2837 DVDD.n103 DVSS 0.051683f
C2838 DVDD.n104 DVSS 0.153995f
C2839 DVDD.n105 DVSS 0.014242f
C2840 DVDD.n106 DVSS 0.027444f
C2841 DVDD.n107 DVSS 0.051683f
C2842 DVDD.n108 DVSS 0.153995f
C2843 DVDD.n109 DVSS 0.014242f
C2844 DVDD.n110 DVSS 0.027444f
C2845 DVDD.n111 DVSS 0.051683f
C2846 DVDD.n112 DVSS 0.153995f
C2847 DVDD.n113 DVSS 0.014242f
C2848 DVDD.n114 DVSS 0.027444f
C2849 DVDD.n115 DVSS 0.051683f
C2850 DVDD.n116 DVSS 0.153995f
C2851 DVDD.n117 DVSS 0.014242f
C2852 DVDD.n118 DVSS 0.027444f
C2853 DVDD.n119 DVSS 0.051683f
C2854 DVDD.n120 DVSS 0.153995f
C2855 VOUT.t31 DVSS 0.155449f
C2856 VOUT.t32 DVSS 0.155449f
C2857 VOUT.n0 DVSS 0.499917f
C2858 VOUT.t30 DVSS 0.155449f
C2859 VOUT.t33 DVSS 0.155449f
C2860 VOUT.n1 DVSS 0.493571f
C2861 VOUT.n2 DVSS 1.43512f
C2862 VOUT.t29 DVSS 0.056979f
C2863 VOUT.t34 DVSS 0.058544f
C2864 VOUT.t18 DVSS 0.056969f
C2865 VOUT.n3 DVSS 1.04422f
C2866 VOUT.t19 DVSS 0.056969f
C2867 VOUT.n4 DVSS 0.557341f
C2868 VOUT.t36 DVSS 0.056969f
C2869 VOUT.n5 DVSS 0.557341f
C2870 VOUT.t13 DVSS 0.056969f
C2871 VOUT.n6 DVSS 0.557341f
C2872 VOUT.t20 DVSS 0.056969f
C2873 VOUT.n7 DVSS 0.557341f
C2874 VOUT.t27 DVSS 0.056969f
C2875 VOUT.n8 DVSS 0.557341f
C2876 VOUT.t9 DVSS 0.056969f
C2877 VOUT.n9 DVSS 0.557341f
C2878 VOUT.t21 DVSS 0.056969f
C2879 VOUT.n10 DVSS 0.557341f
C2880 VOUT.t22 DVSS 0.056969f
C2881 VOUT.n11 DVSS 0.557341f
C2882 VOUT.t24 DVSS 0.056969f
C2883 VOUT.n12 DVSS 0.479543f
C2884 VOUT.t5 DVSS 0.056969f
C2885 VOUT.n13 DVSS 0.709907f
C2886 VOUT.t14 DVSS 0.056969f
C2887 VOUT.n14 DVSS 0.968297f
C2888 VOUT.t23 DVSS 0.056969f
C2889 VOUT.n15 DVSS 0.7937f
C2890 VOUT.t4 DVSS 0.056969f
C2891 VOUT.n16 DVSS 0.829332f
C2892 VOUT.t1 DVSS 0.056969f
C2893 VOUT.n17 DVSS 0.829332f
C2894 VOUT.t26 DVSS 0.056969f
C2895 VOUT.n18 DVSS 0.557341f
C2896 VOUT.t16 DVSS 0.056969f
C2897 VOUT.n19 DVSS 0.557341f
C2898 VOUT.t8 DVSS 0.056969f
C2899 VOUT.n20 DVSS 0.864964f
C2900 VOUT.t0 DVSS 0.056969f
C2901 VOUT.n21 DVSS 0.864964f
C2902 VOUT.t37 DVSS 0.056969f
C2903 VOUT.n22 DVSS 0.557341f
C2904 VOUT.t28 DVSS 0.056969f
C2905 VOUT.n23 DVSS 0.557341f
C2906 VOUT.t12 DVSS 0.056969f
C2907 VOUT.n24 DVSS 0.557341f
C2908 VOUT.t35 DVSS 0.056969f
C2909 VOUT.n25 DVSS 0.557341f
C2910 VOUT.t10 DVSS 0.056969f
C2911 VOUT.n26 DVSS 0.557341f
C2912 VOUT.t17 DVSS 0.056969f
C2913 VOUT.n27 DVSS 0.557341f
C2914 VOUT.t11 DVSS 0.056969f
C2915 VOUT.n28 DVSS 0.810328f
C2916 VOUT.t15 DVSS 0.056969f
C2917 VOUT.n29 DVSS 0.810328f
C2918 VOUT.t3 DVSS 0.056969f
C2919 VOUT.n30 DVSS 0.557341f
C2920 VOUT.t2 DVSS 0.056969f
C2921 VOUT.n31 DVSS 0.557341f
C2922 VOUT.t25 DVSS 0.056969f
C2923 VOUT.n32 DVSS 0.557341f
C2924 VOUT.t7 DVSS 0.056969f
C2925 VOUT.n33 DVSS 0.496171f
C2926 VOUT.n34 DVSS 0.503596f
C2927 VOUT.n35 DVSS 1.62554f
C2928 VOUT.t6 DVSS 0.543589f
C2929 VOUT.n36 DVSS 2.5508f
C2930 VOUT.n37 DVSS 1.07209f
C2931 VOUT.n38 DVSS 1.0633f
C2932 a_16951_764.n0 DVSS 4.89125f
C2933 a_16951_764.n1 DVSS 1.07625f
C2934 a_16951_764.n2 DVSS 4.9015f
C2935 a_16951_764.t2 DVSS 0.176223f
C2936 a_16951_764.t7 DVSS 1.83119f
C2937 a_16951_764.n3 DVSS 0.439579f
C2938 a_16951_764.t4 DVSS 1.83119f
C2939 a_16951_764.n4 DVSS 0.014717f
C2940 a_16951_764.t6 DVSS 1.83119f
C2941 a_16951_764.n5 DVSS 0.015442f
C2942 a_16951_764.t5 DVSS 1.83119f
C2943 a_16951_764.n6 DVSS 1.42285f
C2944 a_16951_764.n7 DVSS 0.978039f
C2945 a_16951_764.t1 DVSS 9.75699f
C2946 a_16951_764.n8 DVSS 0.792274f
C2947 a_16951_764.t3 DVSS 1.52516f
C2948 a_16951_764.n9 DVSS 1.34937f
C2949 a_16951_764.n10 DVSS 0.359396f
C2950 a_16951_764.t0 DVSS 0.176223f
C2951 a_16261_n9984.t21 DVSS 0.228239f
C2952 a_16261_n9984.t16 DVSS 0.051557f
C2953 a_16261_n9984.t23 DVSS 0.051557f
C2954 a_16261_n9984.n0 DVSS 0.148884f
C2955 a_16261_n9984.n1 DVSS 0.534934f
C2956 a_16261_n9984.t14 DVSS 0.051557f
C2957 a_16261_n9984.t17 DVSS 0.051557f
C2958 a_16261_n9984.n2 DVSS 0.148884f
C2959 a_16261_n9984.n3 DVSS 0.291952f
C2960 a_16261_n9984.t25 DVSS 0.051557f
C2961 a_16261_n9984.t24 DVSS 0.051557f
C2962 a_16261_n9984.n4 DVSS 0.148884f
C2963 a_16261_n9984.n5 DVSS 0.291952f
C2964 a_16261_n9984.t19 DVSS 0.051557f
C2965 a_16261_n9984.t18 DVSS 0.051557f
C2966 a_16261_n9984.n6 DVSS 0.148884f
C2967 a_16261_n9984.n7 DVSS 0.291952f
C2968 a_16261_n9984.t27 DVSS 0.051557f
C2969 a_16261_n9984.t15 DVSS 0.051557f
C2970 a_16261_n9984.n8 DVSS 0.148884f
C2971 a_16261_n9984.n9 DVSS 0.292114f
C2972 a_16261_n9984.t20 DVSS 0.051557f
C2973 a_16261_n9984.t26 DVSS 0.051557f
C2974 a_16261_n9984.n10 DVSS 0.148884f
C2975 a_16261_n9984.n11 DVSS 0.389132f
C2976 a_16261_n9984.t22 DVSS 0.180297f
C2977 a_16261_n9984.n12 DVSS 0.545326f
C2978 a_16261_n9984.t8 DVSS 0.081756f
C2979 a_16261_n9984.n13 DVSS 1.13233f
C2980 a_16261_n9984.t5 DVSS 0.081756f
C2981 a_16261_n9984.n14 DVSS 0.799941f
C2982 a_16261_n9984.t10 DVSS 0.084f
C2983 a_16261_n9984.t7 DVSS 0.081756f
C2984 a_16261_n9984.n15 DVSS 1.50022f
C2985 a_16261_n9984.t4 DVSS 0.081756f
C2986 a_16261_n9984.n16 DVSS 0.799941f
C2987 a_16261_n9984.t12 DVSS 0.081756f
C2988 a_16261_n9984.n17 DVSS 0.799941f
C2989 a_16261_n9984.t6 DVSS 0.081756f
C2990 a_16261_n9984.n18 DVSS 0.799941f
C2991 a_16261_n9984.t3 DVSS 0.081756f
C2992 a_16261_n9984.n19 DVSS 0.799941f
C2993 a_16261_n9984.t1 DVSS 0.081756f
C2994 a_16261_n9984.n20 DVSS 0.799941f
C2995 a_16261_n9984.t28 DVSS 0.081756f
C2996 a_16261_n9984.n21 DVSS 0.799941f
C2997 a_16261_n9984.t9 DVSS 0.081756f
C2998 a_16261_n9984.n22 DVSS 0.799941f
C2999 a_16261_n9984.t2 DVSS 0.081756f
C3000 a_16261_n9984.n23 DVSS 0.799941f
C3001 a_16261_n9984.t13 DVSS 0.081756f
C3002 a_16261_n9984.n24 DVSS 0.799941f
C3003 a_16261_n9984.t11 DVSS 0.081756f
C3004 a_16261_n9984.n25 DVSS 0.799941f
C3005 a_16261_n9984.t29 DVSS 0.081756f
C3006 a_16261_n9984.n26 DVSS 0.799941f
C3007 a_16261_n9984.n27 DVSS 0.519464f
C3008 a_16261_n9984.t0 DVSS 0.362233f
C3009 D93v3.n0 DVSS 15.975301f
C3010 D93v3.n1 DVSS 11.1782f
C3011 D93v3.n2 DVSS 9.93091f
C3012 D93v3.n3 DVSS 6.8945f
C3013 D93v3.t0 DVSS 0.037504f
C3014 D93v3.t15 DVSS 0.795146f
C3015 D93v3.t14 DVSS 0.851454f
C3016 D93v3.t17 DVSS 0.847031f
C3017 D93v3.t5 DVSS 0.847031f
C3018 D93v3.t3 DVSS 0.847031f
C3019 D93v3.t27 DVSS 0.847031f
C3020 D93v3.t19 DVSS 0.847031f
C3021 D93v3.t21 DVSS 0.847031f
C3022 D93v3.t7 DVSS 0.847031f
C3023 D93v3.t9 DVSS 0.847031f
C3024 D93v3.t29 DVSS 0.847031f
C3025 D93v3.t23 DVSS 0.847031f
C3026 D93v3.t25 DVSS 0.847031f
C3027 D93v3.t11 DVSS 0.847031f
C3028 D93v3.n4 DVSS 1.39399f
C3029 D93v3.t12 DVSS 0.851454f
C3030 D93v3.t16 DVSS 0.847031f
C3031 D93v3.t4 DVSS 0.847031f
C3032 D93v3.t2 DVSS 0.847031f
C3033 D93v3.t26 DVSS 0.847031f
C3034 D93v3.t18 DVSS 0.847031f
C3035 D93v3.t20 DVSS 0.847031f
C3036 D93v3.t6 DVSS 0.847031f
C3037 D93v3.t8 DVSS 0.847031f
C3038 D93v3.t28 DVSS 0.847031f
C3039 D93v3.t22 DVSS 0.847031f
C3040 D93v3.t24 DVSS 0.847031f
C3041 D93v3.t10 DVSS 0.847031f
C3042 D93v3.t13 DVSS 0.847031f
C3043 D93v3.n5 DVSS 0.031631f
C3044 D93v3.t1 DVSS 0.035219f
C3045 D93v3.n6 DVSS 0.031067f
C3046 ia_opamp_0.V2.t13 DVSS 0.053792f
C3047 ia_opamp_0.V2.t6 DVSS 0.052345f
C3048 ia_opamp_0.V2.n0 DVSS 0.959458f
C3049 ia_opamp_0.V2.t0 DVSS 0.052348f
C3050 ia_opamp_0.V2.n1 DVSS 0.512098f
C3051 ia_opamp_0.V2.t32 DVSS 0.052345f
C3052 ia_opamp_0.V2.n2 DVSS 0.512101f
C3053 ia_opamp_0.V2.t21 DVSS 0.052345f
C3054 ia_opamp_0.V2.n3 DVSS 0.512101f
C3055 ia_opamp_0.V2.t23 DVSS 0.052345f
C3056 ia_opamp_0.V2.n4 DVSS 0.512101f
C3057 ia_opamp_0.V2.t2 DVSS 0.052345f
C3058 ia_opamp_0.V2.n5 DVSS 0.512101f
C3059 ia_opamp_0.V2.t14 DVSS 0.052345f
C3060 ia_opamp_0.V2.n6 DVSS 0.512101f
C3061 ia_opamp_0.V2.t29 DVSS 0.052345f
C3062 ia_opamp_0.V2.n7 DVSS 0.512101f
C3063 ia_opamp_0.V2.t1 DVSS 0.052345f
C3064 ia_opamp_0.V2.n8 DVSS 0.512101f
C3065 ia_opamp_0.V2.t3 DVSS 0.052345f
C3066 ia_opamp_0.V2.n9 DVSS 0.512101f
C3067 ia_opamp_0.V2.t7 DVSS 0.052345f
C3068 ia_opamp_0.V2.n10 DVSS 0.512101f
C3069 ia_opamp_0.V2.t22 DVSS 0.052345f
C3070 ia_opamp_0.V2.n11 DVSS 0.512101f
C3071 ia_opamp_0.V2.t4 DVSS 0.052345f
C3072 ia_opamp_0.V2.n12 DVSS 0.512101f
C3073 ia_opamp_0.V2.t8 DVSS 0.052345f
C3074 ia_opamp_0.V2.n13 DVSS 0.512101f
C3075 ia_opamp_0.V2.t17 DVSS 0.052345f
C3076 ia_opamp_0.V2.n14 DVSS 0.744553f
C3077 ia_opamp_0.V2.t30 DVSS 0.052345f
C3078 ia_opamp_0.V2.n15 DVSS 0.744553f
C3079 ia_opamp_0.V2.t16 DVSS 0.052345f
C3080 ia_opamp_0.V2.n16 DVSS 0.512101f
C3081 ia_opamp_0.V2.t19 DVSS 0.052345f
C3082 ia_opamp_0.V2.n17 DVSS 0.512101f
C3083 ia_opamp_0.V2.t27 DVSS 0.052345f
C3084 ia_opamp_0.V2.n18 DVSS 0.512101f
C3085 ia_opamp_0.V2.t18 DVSS 0.052345f
C3086 ia_opamp_0.V2.n19 DVSS 0.512101f
C3087 ia_opamp_0.V2.t24 DVSS 0.052345f
C3088 ia_opamp_0.V2.n20 DVSS 0.512101f
C3089 ia_opamp_0.V2.t20 DVSS 0.052345f
C3090 ia_opamp_0.V2.n21 DVSS 0.512101f
C3091 ia_opamp_0.V2.t10 DVSS 0.052345f
C3092 ia_opamp_0.V2.n22 DVSS 0.794754f
C3093 ia_opamp_0.V2.t9 DVSS 0.052345f
C3094 ia_opamp_0.V2.n23 DVSS 0.794754f
C3095 ia_opamp_0.V2.t5 DVSS 0.052345f
C3096 ia_opamp_0.V2.n24 DVSS 0.512101f
C3097 ia_opamp_0.V2.t31 DVSS 0.052345f
C3098 ia_opamp_0.V2.n25 DVSS 0.512101f
C3099 ia_opamp_0.V2.t26 DVSS 0.052345f
C3100 ia_opamp_0.V2.n26 DVSS 0.762014f
C3101 ia_opamp_0.V2.t15 DVSS 0.052345f
C3102 ia_opamp_0.V2.n27 DVSS 0.762014f
C3103 ia_opamp_0.V2.t25 DVSS 0.052345f
C3104 ia_opamp_0.V2.n28 DVSS 0.729274f
C3105 ia_opamp_0.V2.t28 DVSS 0.052345f
C3106 ia_opamp_0.V2.n29 DVSS 0.889699f
C3107 ia_opamp_0.V2.t33 DVSS 0.052345f
C3108 ia_opamp_0.V2.n30 DVSS 0.545385f
C3109 ia_opamp_0.V2.t35 DVSS 0.142831f
C3110 ia_opamp_0.V2.t36 DVSS 0.142831f
C3111 ia_opamp_0.V2.n31 DVSS 0.459338f
C3112 ia_opamp_0.V2.t34 DVSS 0.142831f
C3113 ia_opamp_0.V2.t37 DVSS 0.142831f
C3114 ia_opamp_0.V2.n32 DVSS 0.453507f
C3115 ia_opamp_0.V2.n33 DVSS 1.31863f
C3116 ia_opamp_0.V2.n34 DVSS 0.8293f
C3117 ia_opamp_0.V2.t38 DVSS 1.35988f
C3118 ia_opamp_0.V2.n35 DVSS 0.581694f
C3119 ia_opamp_0.V2.n36 DVSS 0.388897f
C3120 ia_opamp_0.V2.n37 DVSS 1.23069f
C3121 ia_opamp_0.V2.t12 DVSS 0.302102f
C3122 ia_opamp_0.V2.t11 DVSS 0.499465f
C3123 ia_opamp_0.V2.n38 DVSS 1.11384f
C3124 ia_opamp_0.V2.n39 DVSS 3.5343f
C3125 ia_opamp_0.V2.n40 DVSS 4.52698f
C3126 VDD.n0 DVSS 1.57578f
C3127 VDD.n1 DVSS 7.17987f
C3128 VDD.n2 DVSS 1.20711f
C3129 VDD.n3 DVSS 1.79361f
C3130 VDD.n4 DVSS 0.483749f
C3131 VDD.n5 DVSS 7.39733f
C3132 VDD.t173 DVSS 5.9327f
C3133 VDD.t171 DVSS 6.38856f
C3134 VDD.n6 DVSS 0.483749f
C3135 VDD.n7 DVSS -4.31569f
C3136 VDD.t18 DVSS 1.08879f
C3137 VDD.t174 DVSS 1.08879f
C3138 VDD.n8 DVSS 3.18938f
C3139 VDD.t163 DVSS 5.93283f
C3140 VDD.n9 DVSS 0.493096f
C3141 VDD.n10 DVSS 0.815382f
C3142 VDD.t231 DVSS 1.37855f
C3143 VDD.n11 DVSS 3.22555f
C3144 VDD.n12 DVSS 1.09327f
C3145 VDD.n13 DVSS 1.09327f
C3146 VDD.t232 DVSS 5.85716f
C3147 VDD.n14 DVSS 2.80605f
C3148 VDD.n15 DVSS 0.685918f
C3149 VDD.n16 DVSS 6.11902f
C3150 VDD.n17 DVSS 5.48804f
C3151 VDD.t227 DVSS 1.37855f
C3152 VDD.t91 DVSS 1.08879f
C3153 VDD.n18 DVSS 3.07752f
C3154 VDD.n19 DVSS 0.493096f
C3155 VDD.n20 DVSS 0.493096f
C3156 VDD.n21 DVSS 1.81902f
C3157 VDD.n22 DVSS -0.487729f
C3158 VDD.n23 DVSS 0.483749f
C3159 VDD.n24 DVSS 0.483749f
C3160 VDD.n25 DVSS 0.973186f
C3161 VDD.t122 DVSS 1.08879f
C3162 VDD.n26 DVSS 0.078954f
C3163 VDD.n27 DVSS 1.79361f
C3164 VDD.n28 DVSS 5.85667f
C3165 VDD.n29 DVSS 0.685918f
C3166 VDD.n30 DVSS 0.165537f
C3167 VDD.n31 DVSS 0.815382f
C3168 VDD.n32 DVSS 5.00963f
C3169 VDD.t23 DVSS 5.93283f
C3170 VDD.t121 DVSS 5.88743f
C3171 VDD.t22 DVSS 1.37855f
C3172 VDD.n33 DVSS 0.864583f
C3173 VDD.n34 DVSS 1.10537f
C3174 VDD.n35 DVSS 1.10537f
C3175 VDD.n36 DVSS 6.94529f
C3176 VDD.n37 DVSS 0.267253f
C3177 VDD.t71 DVSS 1.37855f
C3178 VDD.t73 DVSS 0.379489f
C3179 VDD.t20 DVSS 0.379489f
C3180 VDD.n38 DVSS 1.40778f
C3181 VDD.n39 DVSS 3.69157f
C3182 VDD.n40 DVSS 7.17987f
C3183 VDD.n41 DVSS 0.257963f
C3184 VDD.n42 DVSS 2.69567f
C3185 VDD.n43 DVSS 1.04624f
C3186 VDD.n44 DVSS 0.325883f
C3187 VDD.n45 DVSS 1.79361f
C3188 VDD.n46 DVSS 0.483749f
C3189 VDD.n47 DVSS 0.815382f
C3190 VDD.t47 DVSS 5.93f
C3191 VDD.t49 DVSS 5.93149f
C3192 VDD.n48 DVSS 0.483749f
C3193 VDD.n49 DVSS 0.306781f
C3194 VDD.n50 DVSS -3.47194f
C3195 VDD.t183 DVSS 1.08879f
C3196 VDD.t48 DVSS 1.08879f
C3197 VDD.n51 DVSS 3.18938f
C3198 VDD.t60 DVSS 5.93149f
C3199 VDD.n52 DVSS 0.493096f
C3200 VDD.n53 DVSS 0.815382f
C3201 VDD.t146 DVSS 1.37855f
C3202 VDD.n54 DVSS 0.685918f
C3203 VDD.n55 DVSS 0.864583f
C3204 VDD.n56 DVSS 1.10537f
C3205 VDD.n57 DVSS 1.10537f
C3206 VDD.n58 DVSS 6.94529f
C3207 VDD.n59 DVSS 5.48804f
C3208 VDD.t144 DVSS 1.37855f
C3209 VDD.n60 DVSS 0.809448f
C3210 VDD.t26 DVSS 0.379489f
C3211 VDD.t28 DVSS 0.379489f
C3212 VDD.n61 DVSS 1.40778f
C3213 VDD.n62 DVSS 3.69157f
C3214 VDD.n63 DVSS 4.57059f
C3215 VDD.n64 DVSS 1.79361f
C3216 VDD.n65 DVSS 0.483749f
C3217 VDD.n66 DVSS 0.815382f
C3218 VDD.t111 DVSS 5.93f
C3219 VDD.t29 DVSS 5.93149f
C3220 VDD.n67 DVSS 0.654319f
C3221 VDD.n68 DVSS 0.815382f
C3222 VDD.n69 DVSS 5.1712f
C3223 VDD.t15 DVSS 5.93149f
C3224 VDD.n70 DVSS 0.493096f
C3225 VDD.n71 DVSS 4.00249f
C3226 VDD.n72 DVSS 2.89657f
C3227 VDD.t67 DVSS 1.08879f
C3228 VDD.n73 DVSS 5.85667f
C3229 VDD.n74 DVSS 0.685918f
C3230 VDD.n75 DVSS 2.80492f
C3231 VDD.n76 DVSS 1.09327f
C3232 VDD.n77 DVSS 1.09327f
C3233 VDD.t149 DVSS 5.85583f
C3234 VDD.n78 DVSS 5.79531f
C3235 VDD.n79 DVSS 5.79531f
C3236 VDD.t119 DVSS 7.88343f
C3237 VDD.t147 DVSS 5.85583f
C3238 VDD.n80 DVSS 0.311392f
C3239 VDD.n81 DVSS 0.973186f
C3240 VDD.t118 DVSS 1.37855f
C3241 VDD.n82 DVSS 3.93048f
C3242 VDD.n83 DVSS 0.483749f
C3243 VDD.n84 DVSS 0.815382f
C3244 VDD.t58 DVSS 5.93f
C3245 VDD.n85 DVSS 0.483749f
C3246 VDD.t52 DVSS 1.08879f
C3247 VDD.t59 DVSS 1.08879f
C3248 VDD.n86 DVSS 3.18938f
C3249 VDD.n87 DVSS 2.593f
C3250 VDD.n88 DVSS 0.815382f
C3251 VDD.t135 DVSS 5.93149f
C3252 VDD.t51 DVSS 5.88609f
C3253 VDD.n89 DVSS 1.09327f
C3254 VDD.t178 DVSS 1.37855f
C3255 VDD.n90 DVSS 0.685918f
C3256 VDD.t168 DVSS 0.379489f
C3257 VDD.t176 DVSS 0.379489f
C3258 VDD.n91 DVSS 1.40778f
C3259 VDD.n92 DVSS 3.69157f
C3260 VDD.n93 DVSS 4.57059f
C3261 VDD.n94 DVSS 5.48804f
C3262 VDD.t170 DVSS 1.37855f
C3263 VDD.n95 DVSS 0.809448f
C3264 VDD.n96 DVSS 1.10537f
C3265 VDD.n97 DVSS 1.10537f
C3266 VDD.t4 DVSS 5.93149f
C3267 VDD.n98 DVSS 0.493096f
C3268 VDD.n99 DVSS 0.483749f
C3269 VDD.t5 DVSS 1.08879f
C3270 VDD.n100 DVSS 3.07752f
C3271 VDD.n101 DVSS 0.159917f
C3272 VDD.n102 DVSS 2.80492f
C3273 VDD.n103 DVSS 0.078966f
C3274 VDD.n104 DVSS -0.488632f
C3275 VDD.n105 DVSS 0.483749f
C3276 VDD.n106 DVSS 0.973186f
C3277 VDD.t3 DVSS 1.08879f
C3278 VDD.n107 DVSS 1.79361f
C3279 VDD.n108 DVSS 5.85667f
C3280 VDD.n109 DVSS 0.685918f
C3281 VDD.n110 DVSS 0.559325f
C3282 VDD.n111 DVSS 0.815382f
C3283 VDD.t43 DVSS 5.93149f
C3284 VDD.t2 DVSS 5.88609f
C3285 VDD.t63 DVSS 1.37855f
C3286 VDD.n112 DVSS 0.864583f
C3287 VDD.n113 DVSS 1.10537f
C3288 VDD.n114 DVSS 1.10537f
C3289 VDD.n115 DVSS 2.89657f
C3290 VDD.n116 DVSS 0.704833f
C3291 VDD.t83 DVSS 1.37855f
C3292 VDD.t34 DVSS 0.379489f
C3293 VDD.t65 DVSS 0.379489f
C3294 VDD.n117 DVSS 1.40778f
C3295 VDD.n118 DVSS 3.69157f
C3296 VDD.n119 DVSS 23.788101f
C3297 VDD.n120 DVSS 17.9816f
C3298 VDD.n121 DVSS 11.164001f
C3299 VDD.t246 DVSS 1.06362f
C3300 VDD.t241 DVSS 1.06364f
C3301 VDD.n122 DVSS 8.907041f
C3302 VDD.t247 DVSS 1.06361f
C3303 VDD.t242 DVSS 1.06364f
C3304 VDD.n123 DVSS 8.90681f
C3305 VDD.n124 DVSS 12.372001f
C3306 VDD.n125 DVSS 9.04217f
C3307 VDD.n126 DVSS 12.2864f
C3308 VDD.n127 DVSS 18.333f
C3309 VDD.n128 DVSS 11.8858f
C3310 VDD.n129 DVSS 13.2969f
C3311 VDD.n130 DVSS 13.2969f
C3312 VDD.n131 DVSS 56.4963f
C3313 VDD.n132 DVSS 12.246401f
C3314 VDD.n133 DVSS 11.9066f
C3315 VDD.n134 DVSS 12.3962f
C3316 VDD.n135 DVSS 13.3042f
C3317 VDD.n136 DVSS 56.6275f
C3318 VDD.n137 DVSS 56.4963f
C3319 VDD.n138 DVSS 56.6275f
C3320 VDD.n139 DVSS 13.3042f
C3321 VDD.n140 DVSS 12.3796f
C3322 VDD.n141 DVSS 12.2295f
C3323 VDD.n142 DVSS 11.1439f
C3324 VDD.n143 DVSS 11.677501f
C3325 VDD.n144 DVSS 16.731699f
C3326 VDD.n145 DVSS 6.4881f
C3327 VDD.n146 DVSS 8.74987f
C3328 VDD.n147 DVSS 0.856518f
C3329 VDD.n148 DVSS 3.98477f
C3330 VDD.n149 DVSS 7.595201f
C3331 VDD.t82 DVSS 8.236f
C3332 VDD.t33 DVSS 5.85583f
C3333 VDD.n150 DVSS 3.90389f
C3334 VDD.t64 DVSS 5.85583f
C3335 VDD.t62 DVSS 7.88343f
C3336 VDD.n151 DVSS 5.79531f
C3337 VDD.n152 DVSS 5.79531f
C3338 VDD.n153 DVSS 1.09327f
C3339 VDD.n154 DVSS 3.22555f
C3340 VDD.n155 DVSS -3.47194f
C3341 VDD.n156 DVSS 5.1712f
C3342 VDD.n157 DVSS 0.493096f
C3343 VDD.n158 DVSS 3.90389f
C3344 VDD.n159 DVSS 0.493096f
C3345 VDD.n160 DVSS 0.067995f
C3346 VDD.n161 DVSS 2.593f
C3347 VDD.t44 DVSS 1.08879f
C3348 VDD.n162 DVSS 2.49111f
C3349 VDD.n163 DVSS 4.2323f
C3350 VDD.n164 DVSS 7.17987f
C3351 VDD.t7 DVSS 1.08879f
C3352 VDD.n165 DVSS 3.18938f
C3353 VDD.n166 DVSS 2.26344f
C3354 VDD.n167 DVSS 0.654319f
C3355 VDD.n168 DVSS 4.00249f
C3356 VDD.t6 DVSS 5.93f
C3357 VDD.n169 DVSS 3.90389f
C3358 VDD.n170 DVSS 0.493096f
C3359 VDD.n171 DVSS 0.815382f
C3360 VDD.n172 DVSS 6.94529f
C3361 VDD.n173 DVSS 5.79531f
C3362 VDD.n174 DVSS 5.79531f
C3363 VDD.t177 DVSS 7.88343f
C3364 VDD.t175 DVSS 5.85583f
C3365 VDD.n175 DVSS 3.90389f
C3366 VDD.t167 DVSS 5.85583f
C3367 VDD.t169 DVSS 7.88343f
C3368 VDD.n176 DVSS 6.94529f
C3369 VDD.n177 DVSS 1.09327f
C3370 VDD.n178 DVSS 3.93048f
C3371 VDD.n179 DVSS 0.856518f
C3372 VDD.n180 DVSS 6.11902f
C3373 VDD.t120 DVSS 1.37855f
C3374 VDD.n181 DVSS 3.22555f
C3375 VDD.n182 DVSS 0.864583f
C3376 VDD.t150 DVSS 0.379489f
C3377 VDD.t148 DVSS 0.379489f
C3378 VDD.n183 DVSS 1.40778f
C3379 VDD.n184 DVSS 3.69157f
C3380 VDD.n185 DVSS 0.856518f
C3381 VDD.n186 DVSS 6.11902f
C3382 VDD.n187 DVSS 0.809448f
C3383 VDD.t134 DVSS 1.08879f
C3384 VDD.n188 DVSS 3.07752f
C3385 VDD.n189 DVSS 4.57059f
C3386 VDD.n190 DVSS 7.17987f
C3387 VDD.t136 DVSS 1.08879f
C3388 VDD.n191 DVSS 2.49111f
C3389 VDD.n192 DVSS 4.2323f
C3390 VDD.n193 DVSS 5.85667f
C3391 VDD.n194 DVSS 0.864583f
C3392 VDD.n195 DVSS 3.22555f
C3393 VDD.n196 DVSS 2.26344f
C3394 VDD.n197 DVSS 0.654319f
C3395 VDD.n198 DVSS 4.00249f
C3396 VDD.n199 DVSS -0.488632f
C3397 VDD.n200 DVSS -3.47194f
C3398 VDD.n201 DVSS 5.1712f
C3399 VDD.n202 DVSS 0.493096f
C3400 VDD.n203 DVSS 3.90389f
C3401 VDD.n204 DVSS 0.493096f
C3402 VDD.n205 DVSS 0.067995f
C3403 VDD.n206 DVSS 1.79361f
C3404 VDD.n207 DVSS 0.078966f
C3405 VDD.n208 DVSS 0.493096f
C3406 VDD.t117 DVSS 7.88343f
C3407 VDD.n209 DVSS 6.94529f
C3408 VDD.n210 DVSS 6.94529f
C3409 VDD.t133 DVSS 5.93149f
C3410 VDD.n211 DVSS 3.90389f
C3411 VDD.n212 DVSS 0.493096f
C3412 VDD.n213 DVSS 5.48804f
C3413 VDD.n214 DVSS 2.89657f
C3414 VDD.n215 DVSS 0.311392f
C3415 VDD.n216 DVSS 1.10537f
C3416 VDD.n217 DVSS 3.90389f
C3417 VDD.n218 DVSS 1.10537f
C3418 VDD.n219 DVSS 0.159917f
C3419 VDD.n220 DVSS 0.067995f
C3420 VDD.n221 DVSS 2.593f
C3421 VDD.t16 DVSS 1.08879f
C3422 VDD.n222 DVSS 2.49111f
C3423 VDD.n223 DVSS 4.2323f
C3424 VDD.n224 DVSS 7.17987f
C3425 VDD.t112 DVSS 1.08879f
C3426 VDD.n225 DVSS 3.18938f
C3427 VDD.n226 DVSS 2.26344f
C3428 VDD.n227 DVSS 0.973186f
C3429 VDD.n228 DVSS -3.47194f
C3430 VDD.n229 DVSS -0.488632f
C3431 VDD.t66 DVSS 5.88609f
C3432 VDD.n230 DVSS 3.90389f
C3433 VDD.n231 DVSS 0.493096f
C3434 VDD.n232 DVSS 0.483749f
C3435 VDD.n233 DVSS 0.493096f
C3436 VDD.n234 DVSS 3.90389f
C3437 VDD.n235 DVSS 0.493096f
C3438 VDD.n236 DVSS 0.078966f
C3439 VDD.t30 DVSS 1.08879f
C3440 VDD.n237 DVSS 3.07752f
C3441 VDD.n238 DVSS 2.80492f
C3442 VDD.n239 DVSS 0.159917f
C3443 VDD.n240 DVSS 0.067995f
C3444 VDD.n241 DVSS 2.593f
C3445 VDD.t61 DVSS 1.08879f
C3446 VDD.n242 DVSS 2.49111f
C3447 VDD.n243 DVSS 4.2323f
C3448 VDD.n244 DVSS 5.85667f
C3449 VDD.n245 DVSS 6.11902f
C3450 VDD.n246 DVSS 0.856518f
C3451 VDD.n247 DVSS 3.93048f
C3452 VDD.n248 DVSS 1.09327f
C3453 VDD.n249 DVSS 6.94529f
C3454 VDD.t143 DVSS 7.88343f
C3455 VDD.t25 DVSS 5.85583f
C3456 VDD.n250 DVSS 3.90389f
C3457 VDD.t27 DVSS 5.85583f
C3458 VDD.t145 DVSS 7.88343f
C3459 VDD.n251 DVSS 5.79531f
C3460 VDD.n252 DVSS 5.79531f
C3461 VDD.n253 DVSS 1.09327f
C3462 VDD.n254 DVSS 3.22555f
C3463 VDD.n255 DVSS 5.1712f
C3464 VDD.n256 DVSS 0.493096f
C3465 VDD.n257 DVSS 3.90389f
C3466 VDD.t182 DVSS 5.88609f
C3467 VDD.n258 DVSS -0.488632f
C3468 VDD.n259 DVSS 4.00249f
C3469 VDD.n260 DVSS 0.654319f
C3470 VDD.n261 DVSS 2.26344f
C3471 VDD.n262 DVSS 0.929982f
C3472 VDD.n263 DVSS 2.88865f
C3473 VDD.n264 DVSS 2.89412f
C3474 VDD.n265 DVSS 0.310938f
C3475 VDD.n266 DVSS 0.340093f
C3476 VDD.n267 DVSS 4.37915f
C3477 VDD.n268 DVSS 2.17878f
C3478 VDD.n269 DVSS 0.493096f
C3479 VDD.n270 DVSS 3.90389f
C3480 VDD.n271 DVSS 0.493096f
C3481 VDD.n272 DVSS 0.079072f
C3482 VDD.n273 DVSS 0.263342f
C3483 VDD.n274 DVSS 0.200037f
C3484 VDD.n275 DVSS 0.480165f
C3485 VDD.n276 DVSS 1.36366f
C3486 VDD.t50 DVSS 1.08879f
C3487 VDD.n277 DVSS 1.62913f
C3488 VDD.n278 DVSS 4.57059f
C3489 VDD.n279 DVSS 6.11902f
C3490 VDD.n280 DVSS 0.856518f
C3491 VDD.n281 DVSS 0.916949f
C3492 VDD.n282 DVSS 1.09327f
C3493 VDD.n283 DVSS 6.94529f
C3494 VDD.t70 DVSS 7.88343f
C3495 VDD.t72 DVSS 5.85583f
C3496 VDD.n284 DVSS 3.90389f
C3497 VDD.t19 DVSS 5.85583f
C3498 VDD.t21 DVSS 7.88343f
C3499 VDD.n285 DVSS 4.76637f
C3500 VDD.n286 DVSS 1.09327f
C3501 VDD.n287 DVSS 3.22555f
C3502 VDD.n288 DVSS -3.47194f
C3503 VDD.n289 DVSS 5.1712f
C3504 VDD.n290 DVSS 0.493096f
C3505 VDD.n291 DVSS 3.90477f
C3506 VDD.n292 DVSS 0.493096f
C3507 VDD.n293 DVSS 0.067995f
C3508 VDD.n294 DVSS 2.593f
C3509 VDD.t24 DVSS 1.08879f
C3510 VDD.n295 DVSS 2.49111f
C3511 VDD.n296 DVSS 4.2323f
C3512 VDD.n297 DVSS 4.57059f
C3513 VDD.n298 DVSS 7.17987f
C3514 VDD.t69 DVSS 1.08879f
C3515 VDD.n299 DVSS 3.18938f
C3516 VDD.n300 DVSS 2.26344f
C3517 VDD.n301 DVSS 0.654319f
C3518 VDD.n302 DVSS 0.499445f
C3519 VDD.n303 DVSS 3.98937f
C3520 VDD.t68 DVSS 5.47879f
C3521 VDD.n304 DVSS 3.90477f
C3522 VDD.t90 DVSS 5.93283f
C3523 VDD.t226 DVSS 7.88522f
C3524 VDD.n305 DVSS 6.94686f
C3525 VDD.n306 DVSS 6.94686f
C3526 VDD.n307 DVSS 0.815382f
C3527 VDD.n308 DVSS 0.809448f
C3528 VDD.n309 DVSS 3.93048f
C3529 VDD.n310 DVSS 0.856518f
C3530 VDD.t233 DVSS 0.379489f
C3531 VDD.t229 DVSS 0.379489f
C3532 VDD.n311 DVSS 1.40778f
C3533 VDD.n312 DVSS 3.69157f
C3534 VDD.n313 DVSS 0.864583f
C3535 VDD.n314 DVSS 5.85667f
C3536 VDD.n315 DVSS 4.2323f
C3537 VDD.t164 DVSS 1.08879f
C3538 VDD.n316 DVSS 2.49111f
C3539 VDD.n317 DVSS 0.067995f
C3540 VDD.n318 DVSS 2.593f
C3541 VDD.n319 DVSS 0.159917f
C3542 VDD.n320 DVSS 1.10537f
C3543 VDD.n321 DVSS 5.615f
C3544 VDD.t37 DVSS 4.78702f
C3545 VDD.n322 DVSS 1.35175f
C3546 VDD.t39 DVSS 4.78702f
C3547 VDD.t78 DVSS 6.38269f
C3548 VDD.t76 DVSS 6.38269f
C3549 VDD.t186 DVSS 6.38269f
C3550 VDD.t184 DVSS 6.38269f
C3551 VDD.t137 DVSS 6.73872f
C3552 VDD.n323 DVSS 6.66103f
C3553 VDD.n324 DVSS 6.66103f
C3554 VDD.t138 DVSS 1.22797f
C3555 VDD.t185 DVSS 0.299597f
C3556 VDD.t187 DVSS 0.299597f
C3557 VDD.n325 DVSS 0.746184f
C3558 VDD.t77 DVSS 0.299597f
C3559 VDD.t79 DVSS 0.299597f
C3560 VDD.n326 DVSS 0.746184f
C3561 VDD.t38 DVSS 0.299597f
C3562 VDD.t40 DVSS 0.299597f
C3563 VDD.n327 DVSS 0.746184f
C3564 VDD.t75 DVSS 0.299597f
C3565 VDD.t132 DVSS 0.299597f
C3566 VDD.n328 DVSS 0.746184f
C3567 VDD.t140 DVSS 0.299597f
C3568 VDD.t142 DVSS 0.299597f
C3569 VDD.n329 DVSS 0.746184f
C3570 VDD.t130 DVSS 0.019973f
C3571 VDD.t116 DVSS 0.019973f
C3572 VDD.n330 DVSS 0.045455f
C3573 VDD.t36 DVSS 1.22878f
C3574 VDD.n331 DVSS 3.91367f
C3575 VDD.n332 DVSS 2.90397f
C3576 VDD.n333 DVSS 4.61086f
C3577 VDD.n334 DVSS 5.33543f
C3578 VDD.n335 DVSS 5.33543f
C3579 VDD.n336 DVSS 5.33543f
C3580 VDD.n337 DVSS 5.33543f
C3581 VDD.n338 DVSS 6.3896f
C3582 VDD.n339 DVSS 2.50354f
C3583 VDD.n340 DVSS 0.743567f
C3584 VDD.n341 DVSS 2.67271f
C3585 VDD.n342 DVSS 0.796975f
C3586 VDD.n343 DVSS 2.54985f
C3587 VDD.n344 DVSS 1.26566f
C3588 VDD.n345 DVSS 1.05999f
C3589 VDD.n346 DVSS 1.42195f
C3590 VDD.n347 DVSS 1.42195f
C3591 VDD.t74 DVSS 6.38269f
C3592 VDD.t131 DVSS 6.38269f
C3593 VDD.t139 DVSS 6.38269f
C3594 VDD.t141 DVSS 4.78702f
C3595 VDD.t35 DVSS 5.14305f
C3596 VDD.t129 DVSS 1.16779f
C3597 VDD.t115 DVSS 1.16779f
C3598 VDD.n348 DVSS 0.668392f
C3599 VDD.n349 DVSS 1.05463f
C3600 VDD.n350 DVSS 0.275154f
C3601 VDD.n351 DVSS 3.89678f
C3602 VDD.n352 DVSS 0.275154f
C3603 VDD.n353 DVSS 0.717379f
C3604 VDD.n354 DVSS 0.923181f
C3605 VDD.n355 DVSS 1.93708f
C3606 VDD.n356 DVSS 1.35175f
C3607 VDD.n357 DVSS 5.00752f
C3608 VDD.n358 DVSS 4.16206f
C3609 VDD.t230 DVSS 7.88522f
C3610 VDD.t228 DVSS 5.85716f
C3611 VDD.n359 DVSS 3.90477f
C3612 VDD.n360 DVSS 1.10537f
C3613 VDD.n361 DVSS 0.28555f
C3614 VDD.n362 DVSS 2.83953f
C3615 VDD.n363 DVSS 5.02634f
C3616 VDD.n364 DVSS 0.493096f
C3617 VDD.n365 DVSS 3.90477f
C3618 VDD.t17 DVSS 5.88743f
C3619 VDD.n366 DVSS -0.487729f
C3620 VDD.n367 DVSS 4.01383f
C3621 VDD.n368 DVSS 0.654319f
C3622 VDD.n369 DVSS 2.26344f
C3623 VDD.n370 DVSS 1.87284f
C3624 VDD.n371 DVSS 3.61877f
C3625 VDD.n372 DVSS 0.493096f
C3626 VDD.n373 DVSS 3.90477f
C3627 VDD.n374 DVSS 0.493096f
C3628 VDD.n375 DVSS 0.439662f
C3629 VDD.t172 DVSS 1.08879f
C3630 VDD.n376 DVSS 1.86727f
C3631 VDD.n377 DVSS 6.19271f
C3632 VDD.n378 DVSS 0.02248f
C3633 VDD.n379 DVSS 0.02248f
C3634 VDD.t41 DVSS 2.58294f
C3635 VDD.t152 DVSS 1.05709f
C3636 VDD.n380 DVSS 0.014224f
C3637 VDD.n384 DVSS 0.02248f
C3638 VDD.n385 DVSS 0.02248f
C3639 VDD.n386 DVSS 0.082978f
C3640 VDD.t235 DVSS 0.244327f
C3641 VDD.t203 DVSS 0.067409f
C3642 VDD.n387 DVSS 0.156668f
C3643 VDD.n388 DVSS 0.02248f
C3644 VDD.t151 DVSS 0.038224f
C3645 VDD.t42 DVSS 0.028927f
C3646 VDD.n389 DVSS 0.079201f
C3647 VDD.n390 DVSS 0.013612f
C3648 VDD.n391 DVSS 0.02248f
C3649 VDD.n392 DVSS 0.02248f
C3650 VDD.n393 DVSS 0.02248f
C3651 VDD.n394 DVSS 0.02841f
C3652 VDD.t191 DVSS 0.047825f
C3653 VDD.n395 DVSS 0.059733f
C3654 VDD.n396 DVSS 0.02248f
C3655 VDD.n397 DVSS 0.02248f
C3656 VDD.t31 DVSS 2.58294f
C3657 VDD.t127 DVSS 1.05709f
C3658 VDD.n398 DVSS 0.014224f
C3659 VDD.n402 DVSS 0.02248f
C3660 VDD.n403 DVSS 0.02248f
C3661 VDD.n404 DVSS 0.082647f
C3662 VDD.t248 DVSS 0.244327f
C3663 VDD.t155 DVSS 0.067409f
C3664 VDD.n405 DVSS 0.156668f
C3665 VDD.n406 DVSS 0.02248f
C3666 VDD.t126 DVSS 0.038224f
C3667 VDD.t32 DVSS 0.028927f
C3668 VDD.n407 DVSS 0.079201f
C3669 VDD.n408 DVSS 0.013612f
C3670 VDD.n409 DVSS 0.02248f
C3671 VDD.n410 DVSS 0.02248f
C3672 VDD.n411 DVSS 0.02248f
C3673 VDD.n412 DVSS 0.02841f
C3674 VDD.t46 DVSS 0.047825f
C3675 VDD.n413 DVSS 0.059733f
C3676 VDD.n414 DVSS 0.02248f
C3677 VDD.n415 DVSS 0.02248f
C3678 VDD.t96 DVSS 2.58294f
C3679 VDD.t98 DVSS 1.05709f
C3680 VDD.n416 DVSS 0.014224f
C3681 VDD.n420 DVSS 0.02248f
C3682 VDD.n421 DVSS 0.02248f
C3683 VDD.n422 DVSS 0.082647f
C3684 VDD.t239 DVSS 0.244327f
C3685 VDD.t215 DVSS 0.067409f
C3686 VDD.n423 DVSS 0.156668f
C3687 VDD.n424 DVSS 0.02248f
C3688 VDD.t97 DVSS 0.038224f
C3689 VDD.t165 DVSS 0.028927f
C3690 VDD.n425 DVSS 0.079201f
C3691 VDD.n426 DVSS 0.013612f
C3692 VDD.n427 DVSS 0.02248f
C3693 VDD.n428 DVSS 0.02248f
C3694 VDD.n429 DVSS 0.02248f
C3695 VDD.n430 DVSS 0.02841f
C3696 VDD.t201 DVSS 0.047825f
C3697 VDD.n431 DVSS 0.059733f
C3698 VDD.n432 DVSS 0.02248f
C3699 VDD.n433 DVSS 0.02248f
C3700 VDD.t107 DVSS 2.58294f
C3701 VDD.t193 DVSS 1.05709f
C3702 VDD.n434 DVSS 0.014224f
C3703 VDD.n438 DVSS 0.02248f
C3704 VDD.n439 DVSS 0.02248f
C3705 VDD.n440 DVSS 0.082647f
C3706 VDD.t243 DVSS 0.244327f
C3707 VDD.t221 DVSS 0.067409f
C3708 VDD.n441 DVSS 0.156668f
C3709 VDD.n442 DVSS 0.02248f
C3710 VDD.t192 DVSS 0.038224f
C3711 VDD.t108 DVSS 0.028927f
C3712 VDD.n443 DVSS 0.079201f
C3713 VDD.n444 DVSS 0.013612f
C3714 VDD.n445 DVSS 0.02248f
C3715 VDD.n446 DVSS 0.02248f
C3716 VDD.n447 DVSS 0.02248f
C3717 VDD.n448 DVSS 0.02841f
C3718 VDD.t95 DVSS 0.047825f
C3719 VDD.n449 DVSS 0.059733f
C3720 VDD.n450 DVSS 0.02248f
C3721 VDD.n451 DVSS 0.02248f
C3722 VDD.n452 DVSS 0.015342f
C3723 VDD.n453 DVSS 0.02248f
C3724 VDD.n454 DVSS 0.02248f
C3725 VDD.n455 DVSS 0.082647f
C3726 VDD.t236 DVSS 0.244327f
C3727 VDD.t212 DVSS 0.067409f
C3728 VDD.n456 DVSS 0.156668f
C3729 VDD.n457 DVSS 0.033908f
C3730 VDD.n458 DVSS 0.041324f
C3731 VDD.n459 DVSS 0.062846f
C3732 VDD.n460 DVSS 0.041324f
C3733 VDD.n461 DVSS 0.088433f
C3734 VDD.n462 DVSS 0.170494f
C3735 VDD.t213 DVSS 0.072182f
C3736 VDD.n463 DVSS 0.129401f
C3737 VDD.n464 DVSS 0.041324f
C3738 VDD.n465 DVSS 0.073177f
C3739 VDD.n466 DVSS 0.02248f
C3740 VDD.n467 DVSS 0.02248f
C3741 VDD.t211 DVSS 1.47253f
C3742 VDD.n469 DVSS 2.19935f
C3743 VDD.n470 DVSS 0.022012f
C3744 VDD.n471 DVSS 0.037467f
C3745 VDD.n472 DVSS 0.055959f
C3746 VDD.n473 DVSS 0.025585f
C3747 VDD.n474 DVSS 0.014636f
C3748 VDD.n475 DVSS 1.32039f
C3749 VDD.t194 DVSS 0.028448f
C3750 VDD.n476 DVSS 0.049105f
C3751 VDD.n477 DVSS 0.02358f
C3752 VDD.n478 DVSS 0.034436f
C3753 VDD.n479 DVSS 0.065858f
C3754 VDD.n480 DVSS 0.014636f
C3755 VDD.n481 DVSS 0.068873f
C3756 VDD.n482 DVSS 0.02248f
C3757 VDD.n483 DVSS 0.02248f
C3758 VDD.n484 DVSS 0.02248f
C3759 VDD.n485 DVSS 0.02248f
C3760 VDD.n486 DVSS 0.014636f
C3761 VDD.n487 DVSS 0.068012f
C3762 VDD.n488 DVSS 0.210629f
C3763 VDD.n489 DVSS 0.055959f
C3764 VDD.n490 DVSS 0.026688f
C3765 VDD.n491 DVSS 0.082647f
C3766 VDD.n492 DVSS 0.01686f
C3767 VDD.n493 DVSS 0.02248f
C3768 VDD.n494 DVSS 0.02248f
C3769 VDD.n495 DVSS 0.01686f
C3770 VDD.n496 DVSS 0.082647f
C3771 VDD.n497 DVSS 0.041324f
C3772 VDD.n498 DVSS 0.062846f
C3773 VDD.n499 DVSS 0.041324f
C3774 VDD.n500 DVSS 0.088433f
C3775 VDD.n501 DVSS 0.170494f
C3776 VDD.t222 DVSS 0.072182f
C3777 VDD.n502 DVSS 0.129401f
C3778 VDD.n503 DVSS 0.041324f
C3779 VDD.n504 DVSS 0.073177f
C3780 VDD.n505 DVSS 0.02248f
C3781 VDD.n506 DVSS 0.02248f
C3782 VDD.t94 DVSS 0.687584f
C3783 VDD.t220 DVSS 0.999688f
C3784 VDD.n508 DVSS 1.36799f
C3785 VDD.n509 DVSS 0.022012f
C3786 VDD.n510 DVSS 0.037467f
C3787 VDD.n511 DVSS 0.055959f
C3788 VDD.n512 DVSS 0.025585f
C3789 VDD.n513 DVSS 0.014636f
C3790 VDD.n514 DVSS 1.32039f
C3791 VDD.t99 DVSS 0.028448f
C3792 VDD.n515 DVSS 0.049105f
C3793 VDD.n516 DVSS 0.02358f
C3794 VDD.n517 DVSS 0.034436f
C3795 VDD.n518 DVSS 0.065858f
C3796 VDD.n519 DVSS 0.014636f
C3797 VDD.n520 DVSS 0.068873f
C3798 VDD.n521 DVSS 0.02248f
C3799 VDD.n522 DVSS 0.02248f
C3800 VDD.n523 DVSS 0.02248f
C3801 VDD.n524 DVSS 0.02248f
C3802 VDD.n525 DVSS 0.014636f
C3803 VDD.n526 DVSS 0.068012f
C3804 VDD.n527 DVSS 0.210629f
C3805 VDD.n528 DVSS 0.055959f
C3806 VDD.n529 DVSS 0.026688f
C3807 VDD.n530 DVSS 0.082647f
C3808 VDD.n531 DVSS 0.01686f
C3809 VDD.n532 DVSS 0.02248f
C3810 VDD.n533 DVSS 0.02248f
C3811 VDD.n534 DVSS 0.01686f
C3812 VDD.n535 DVSS 0.082647f
C3813 VDD.n536 DVSS 0.041324f
C3814 VDD.n537 DVSS 0.062846f
C3815 VDD.n538 DVSS 0.041324f
C3816 VDD.n539 DVSS 0.088433f
C3817 VDD.n540 DVSS 0.170494f
C3818 VDD.t216 DVSS 0.072182f
C3819 VDD.n541 DVSS 0.129401f
C3820 VDD.n542 DVSS 0.041324f
C3821 VDD.n543 DVSS 0.073177f
C3822 VDD.n544 DVSS 0.02248f
C3823 VDD.n545 DVSS 0.02248f
C3824 VDD.t200 DVSS 0.687584f
C3825 VDD.t214 DVSS 0.999688f
C3826 VDD.n547 DVSS 1.36799f
C3827 VDD.n548 DVSS 0.022012f
C3828 VDD.n549 DVSS 0.037467f
C3829 VDD.n550 DVSS 0.055959f
C3830 VDD.n551 DVSS 0.025585f
C3831 VDD.n552 DVSS 0.014636f
C3832 VDD.n553 DVSS 1.32039f
C3833 VDD.t128 DVSS 0.028448f
C3834 VDD.n554 DVSS 0.049105f
C3835 VDD.n555 DVSS 0.02358f
C3836 VDD.n556 DVSS 0.034436f
C3837 VDD.n557 DVSS 0.065858f
C3838 VDD.n558 DVSS 0.014636f
C3839 VDD.n559 DVSS 0.068873f
C3840 VDD.n560 DVSS 0.02248f
C3841 VDD.n561 DVSS 0.02248f
C3842 VDD.n562 DVSS 0.02248f
C3843 VDD.n563 DVSS 0.02248f
C3844 VDD.n564 DVSS 0.014636f
C3845 VDD.n565 DVSS 0.068012f
C3846 VDD.n566 DVSS 0.210629f
C3847 VDD.n567 DVSS 0.055959f
C3848 VDD.n568 DVSS 0.026688f
C3849 VDD.n569 DVSS 0.082647f
C3850 VDD.n570 DVSS 0.01686f
C3851 VDD.n571 DVSS 0.02248f
C3852 VDD.n572 DVSS 0.02248f
C3853 VDD.n573 DVSS 0.01686f
C3854 VDD.n574 DVSS 0.082647f
C3855 VDD.n575 DVSS 0.041324f
C3856 VDD.n576 DVSS 0.062846f
C3857 VDD.n577 DVSS 0.041324f
C3858 VDD.n578 DVSS 0.088433f
C3859 VDD.n579 DVSS 0.170494f
C3860 VDD.t156 DVSS 0.072182f
C3861 VDD.n580 DVSS 0.129401f
C3862 VDD.n581 DVSS 0.041324f
C3863 VDD.n582 DVSS 0.073177f
C3864 VDD.n583 DVSS 0.02248f
C3865 VDD.n584 DVSS 0.02248f
C3866 VDD.t45 DVSS 0.687584f
C3867 VDD.t154 DVSS 0.999688f
C3868 VDD.n586 DVSS 1.36799f
C3869 VDD.n587 DVSS 0.022012f
C3870 VDD.n588 DVSS 0.037467f
C3871 VDD.n589 DVSS 0.055959f
C3872 VDD.n590 DVSS 0.025585f
C3873 VDD.n591 DVSS 0.014636f
C3874 VDD.n592 DVSS 1.32039f
C3875 VDD.t153 DVSS 0.028448f
C3876 VDD.n593 DVSS 0.049105f
C3877 VDD.n594 DVSS 0.02358f
C3878 VDD.n595 DVSS 0.034436f
C3879 VDD.n596 DVSS 0.065858f
C3880 VDD.n597 DVSS 0.014636f
C3881 VDD.n598 DVSS 0.068873f
C3882 VDD.n599 DVSS 0.02248f
C3883 VDD.n600 DVSS 0.02248f
C3884 VDD.n601 DVSS 0.02248f
C3885 VDD.n602 DVSS 0.02248f
C3886 VDD.n603 DVSS 0.014636f
C3887 VDD.n604 DVSS 0.068012f
C3888 VDD.n605 DVSS 0.210629f
C3889 VDD.n606 DVSS 0.055959f
C3890 VDD.n607 DVSS 0.026688f
C3891 VDD.n608 DVSS 0.082647f
C3892 VDD.n609 DVSS 0.01686f
C3893 VDD.n610 DVSS 0.02248f
C3894 VDD.n611 DVSS 0.02248f
C3895 VDD.n612 DVSS 0.01686f
C3896 VDD.n613 DVSS 0.082647f
C3897 VDD.n614 DVSS 0.041324f
C3898 VDD.n615 DVSS 0.031854f
C3899 VDD.n616 DVSS 0.07244f
C3900 VDD.n617 DVSS 0.033706f
C3901 VDD.n618 DVSS 0.088433f
C3902 VDD.n619 DVSS 0.170494f
C3903 VDD.t204 DVSS 0.072182f
C3904 VDD.n620 DVSS 0.129401f
C3905 VDD.n621 DVSS 0.041482f
C3906 VDD.n622 DVSS 0.073467f
C3907 VDD.n623 DVSS 0.02248f
C3908 VDD.n624 DVSS 0.02248f
C3909 VDD.t190 DVSS 0.687584f
C3910 VDD.t202 DVSS 0.999688f
C3911 VDD.n626 DVSS 1.36799f
C3912 VDD.n627 DVSS 0.022012f
C3913 VDD.n628 DVSS 0.037467f
C3914 VDD.n629 DVSS 0.05618f
C3915 VDD.n630 DVSS 0.014636f
C3916 VDD.t199 DVSS 0.047825f
C3917 VDD.n631 DVSS 0.059733f
C3918 VDD.n632 DVSS 0.034436f
C3919 VDD.n633 DVSS 0.065858f
C3920 VDD.n634 DVSS 0.014636f
C3921 VDD.n635 DVSS 0.025585f
C3922 VDD.n636 DVSS 0.02248f
C3923 VDD.n637 DVSS 0.02248f
C3924 VDD.n638 DVSS 0.02248f
C3925 VDD.n639 DVSS 0.014636f
C3926 VDD.n640 DVSS 0.02248f
C3927 VDD.n641 DVSS 0.02248f
C3928 VDD.n642 DVSS 0.02248f
C3929 VDD.n643 DVSS 0.02248f
C3930 VDD.n644 DVSS 0.02248f
C3931 VDD.n645 DVSS 0.041324f
C3932 VDD.t161 DVSS 0.067409f
C3933 VDD.n646 DVSS 0.156668f
C3934 VDD.t234 DVSS 0.244327f
C3935 VDD.t162 DVSS 0.072182f
C3936 VDD.n647 DVSS 0.073177f
C3937 VDD.n648 DVSS 0.02248f
C3938 VDD.t102 DVSS 2.58294f
C3939 VDD.t196 DVSS 1.05709f
C3940 VDD.n649 DVSS 0.014224f
C3941 VDD.n650 DVSS 0.02248f
C3942 VDD.n654 DVSS 0.02248f
C3943 VDD.t198 DVSS 0.687584f
C3944 VDD.t160 DVSS 0.999688f
C3945 VDD.n656 DVSS 1.36799f
C3946 VDD.n657 DVSS 0.022012f
C3947 VDD.n658 DVSS 0.014636f
C3948 VDD.t101 DVSS 0.047825f
C3949 VDD.n659 DVSS 0.059733f
C3950 VDD.n660 DVSS 0.034436f
C3951 VDD.n661 DVSS 0.065858f
C3952 VDD.n662 DVSS 0.014636f
C3953 VDD.n663 DVSS 0.025585f
C3954 VDD.n664 DVSS 0.02248f
C3955 VDD.n665 DVSS 0.02248f
C3956 VDD.n666 DVSS 0.02248f
C3957 VDD.n667 DVSS 0.014636f
C3958 VDD.n668 DVSS 0.02248f
C3959 VDD.n669 DVSS 0.02248f
C3960 VDD.n670 DVSS 0.02248f
C3961 VDD.n671 DVSS 0.02248f
C3962 VDD.n672 DVSS 0.02248f
C3963 VDD.n673 DVSS 0.041324f
C3964 VDD.t209 DVSS 0.067409f
C3965 VDD.n674 DVSS 0.156668f
C3966 VDD.t238 DVSS 0.244327f
C3967 VDD.t210 DVSS 0.072182f
C3968 VDD.n675 DVSS 0.073177f
C3969 VDD.n676 DVSS 0.02248f
C3970 VDD.t113 DVSS 2.58294f
C3971 VDD.t179 DVSS 1.05709f
C3972 VDD.n677 DVSS 0.014224f
C3973 VDD.n678 DVSS 0.02248f
C3974 VDD.n682 DVSS 0.02248f
C3975 VDD.t100 DVSS 0.687584f
C3976 VDD.t208 DVSS 0.999688f
C3977 VDD.n684 DVSS 1.36799f
C3978 VDD.n685 DVSS 0.022012f
C3979 VDD.n686 DVSS 0.014636f
C3980 VDD.t54 DVSS 0.047825f
C3981 VDD.n687 DVSS 0.059733f
C3982 VDD.n688 DVSS 0.034436f
C3983 VDD.n689 DVSS 0.065858f
C3984 VDD.n690 DVSS 0.014636f
C3985 VDD.n691 DVSS 0.025585f
C3986 VDD.n692 DVSS 0.02248f
C3987 VDD.n693 DVSS 0.02248f
C3988 VDD.n694 DVSS 0.02248f
C3989 VDD.n695 DVSS 0.014636f
C3990 VDD.n696 DVSS 0.02248f
C3991 VDD.n697 DVSS 0.02248f
C3992 VDD.n698 DVSS 0.02248f
C3993 VDD.n699 DVSS 0.02248f
C3994 VDD.n700 DVSS 0.02248f
C3995 VDD.n701 DVSS 0.041324f
C3996 VDD.t206 DVSS 0.067409f
C3997 VDD.n702 DVSS 0.156668f
C3998 VDD.t237 DVSS 0.244327f
C3999 VDD.t207 DVSS 0.072182f
C4000 VDD.n703 DVSS 0.073177f
C4001 VDD.n704 DVSS 0.02248f
C4002 VDD.t8 DVSS 2.58294f
C4003 VDD.t55 DVSS 1.05709f
C4004 VDD.n705 DVSS 0.014224f
C4005 VDD.n706 DVSS 0.02248f
C4006 VDD.n710 DVSS 0.02248f
C4007 VDD.t53 DVSS 0.687584f
C4008 VDD.t205 DVSS 0.999688f
C4009 VDD.n712 DVSS 1.36799f
C4010 VDD.n713 DVSS 0.022012f
C4011 VDD.n714 DVSS 0.014636f
C4012 VDD.t81 DVSS 0.047825f
C4013 VDD.n715 DVSS 0.059733f
C4014 VDD.n716 DVSS 0.034436f
C4015 VDD.n717 DVSS 0.065858f
C4016 VDD.n718 DVSS 0.014636f
C4017 VDD.n719 DVSS 0.025585f
C4018 VDD.n720 DVSS 0.02248f
C4019 VDD.n721 DVSS 0.02248f
C4020 VDD.n722 DVSS 0.02248f
C4021 VDD.n723 DVSS 0.014636f
C4022 VDD.n724 DVSS 0.02248f
C4023 VDD.n725 DVSS 0.02248f
C4024 VDD.n726 DVSS 0.02248f
C4025 VDD.n727 DVSS 0.02248f
C4026 VDD.n728 DVSS 0.02248f
C4027 VDD.n729 DVSS 0.041324f
C4028 VDD.t158 DVSS 0.067409f
C4029 VDD.n730 DVSS 0.156668f
C4030 VDD.t245 DVSS 0.244327f
C4031 VDD.t159 DVSS 0.072182f
C4032 VDD.n731 DVSS 0.073177f
C4033 VDD.n732 DVSS 0.02248f
C4034 VDD.t88 DVSS 2.58294f
C4035 VDD.t86 DVSS 1.05709f
C4036 VDD.n733 DVSS 0.014224f
C4037 VDD.n734 DVSS 0.02248f
C4038 VDD.n738 DVSS 0.02248f
C4039 VDD.t80 DVSS 0.687584f
C4040 VDD.t157 DVSS 0.999688f
C4041 VDD.n740 DVSS 1.36799f
C4042 VDD.n741 DVSS 0.022012f
C4043 VDD.n742 DVSS 0.014636f
C4044 VDD.t110 DVSS 0.047825f
C4045 VDD.n743 DVSS 0.059733f
C4046 VDD.n744 DVSS 0.034436f
C4047 VDD.n745 DVSS 0.065858f
C4048 VDD.n746 DVSS 0.014636f
C4049 VDD.n747 DVSS 0.025585f
C4050 VDD.n748 DVSS 0.02248f
C4051 VDD.n749 DVSS 0.02248f
C4052 VDD.n750 DVSS 0.02248f
C4053 VDD.n751 DVSS 0.014636f
C4054 VDD.n752 DVSS 0.02248f
C4055 VDD.n753 DVSS 0.02248f
C4056 VDD.n754 DVSS 0.02248f
C4057 VDD.n755 DVSS 0.02248f
C4058 VDD.n756 DVSS 0.02248f
C4059 VDD.n757 DVSS 0.041324f
C4060 VDD.t218 DVSS 0.067409f
C4061 VDD.n758 DVSS 0.156668f
C4062 VDD.t240 DVSS 0.244327f
C4063 VDD.t219 DVSS 0.072182f
C4064 VDD.n759 DVSS 0.073177f
C4065 VDD.n760 DVSS 0.02248f
C4066 VDD.t188 DVSS 2.58294f
C4067 VDD.t223 DVSS 1.05709f
C4068 VDD.n761 DVSS 0.014224f
C4069 VDD.n762 DVSS 0.02248f
C4070 VDD.n766 DVSS 0.02248f
C4071 VDD.t109 DVSS 0.687584f
C4072 VDD.t217 DVSS 0.999688f
C4073 VDD.n768 DVSS 1.36799f
C4074 VDD.n769 DVSS 0.022012f
C4075 VDD.n770 DVSS 0.014636f
C4076 VDD.t93 DVSS 0.047825f
C4077 VDD.n771 DVSS 0.059733f
C4078 VDD.n772 DVSS 0.034436f
C4079 VDD.n773 DVSS 0.065858f
C4080 VDD.n774 DVSS 0.014636f
C4081 VDD.n775 DVSS 0.025585f
C4082 VDD.n776 DVSS 0.02248f
C4083 VDD.n777 DVSS 0.02248f
C4084 VDD.n778 DVSS 0.02248f
C4085 VDD.n779 DVSS 0.014636f
C4086 VDD.n780 DVSS 0.02248f
C4087 VDD.n781 DVSS 0.02248f
C4088 VDD.n782 DVSS 0.02248f
C4089 VDD.n783 DVSS 0.02248f
C4090 VDD.n784 DVSS 0.02248f
C4091 VDD.n785 DVSS 0.041324f
C4092 VDD.t105 DVSS 0.067409f
C4093 VDD.n786 DVSS 0.156668f
C4094 VDD.t244 DVSS 0.244327f
C4095 VDD.t106 DVSS 0.072182f
C4096 VDD.n787 DVSS 0.073177f
C4097 VDD.n788 DVSS 0.02248f
C4098 VDD.t84 DVSS 2.58294f
C4099 VDD.t123 DVSS 1.05709f
C4100 VDD.n789 DVSS 0.014224f
C4101 VDD.n790 DVSS 0.02248f
C4102 VDD.n794 DVSS 0.02248f
C4103 VDD.t92 DVSS 0.687584f
C4104 VDD.t104 DVSS 0.999688f
C4105 VDD.n796 DVSS 1.36799f
C4106 VDD.n797 DVSS 0.022012f
C4107 VDD.n798 DVSS 0.014636f
C4108 VDD.t11 DVSS 0.047825f
C4109 VDD.n799 DVSS 0.059733f
C4110 VDD.n800 DVSS 0.034436f
C4111 VDD.n801 DVSS 0.065858f
C4112 VDD.n802 DVSS 0.014636f
C4113 VDD.n803 DVSS 0.025585f
C4114 VDD.n804 DVSS 0.02248f
C4115 VDD.n805 DVSS 0.02248f
C4116 VDD.n806 DVSS 0.02248f
C4117 VDD.n807 DVSS 0.014636f
C4118 VDD.n808 DVSS 0.02248f
C4119 VDD.t0 DVSS 1.69406f
C4120 VDD.t12 DVSS 0.693308f
C4121 VDD.n809 DVSS 0.014224f
C4122 VDD.n810 DVSS 0.02248f
C4123 VDD.t10 DVSS 1.18422f
C4124 VDD.n812 DVSS 1.01016f
C4125 VDD.n813 DVSS 0.015342f
C4126 VDD.n814 DVSS 0.038713f
C4127 VDD.n815 DVSS 0.082647f
C4128 VDD.n816 DVSS 0.023998f
C4129 VDD.n817 DVSS 0.02248f
C4130 VDD.n818 DVSS 0.026688f
C4131 VDD.n819 DVSS 0.055959f
C4132 VDD.t14 DVSS 0.038224f
C4133 VDD.t1 DVSS 0.028927f
C4134 VDD.n820 DVSS 0.079201f
C4135 VDD.n821 DVSS 0.013612f
C4136 VDD.n822 DVSS 0.210629f
C4137 VDD.n823 DVSS 0.068012f
C4138 VDD.n824 DVSS 0.068873f
C4139 VDD.n825 DVSS 0.02248f
C4140 VDD.n826 DVSS 0.02248f
C4141 VDD.n827 DVSS 0.02841f
C4142 VDD.n828 DVSS 0.02358f
C4143 VDD.t13 DVSS 0.028448f
C4144 VDD.n829 DVSS 0.049105f
C4145 VDD.n830 DVSS 1.32039f
C4146 VDD.n831 DVSS 0.055959f
C4147 VDD.n832 DVSS 0.037467f
C4148 VDD.n833 DVSS 0.02248f
C4149 VDD.n834 DVSS 0.082647f
C4150 VDD.n835 DVSS 0.041324f
C4151 VDD.n836 DVSS 0.129401f
C4152 VDD.n837 DVSS 0.170494f
C4153 VDD.n838 DVSS 0.088433f
C4154 VDD.n839 DVSS 0.041324f
C4155 VDD.n840 DVSS 0.062846f
C4156 VDD.n841 DVSS 0.02248f
C4157 VDD.n842 DVSS 0.01686f
C4158 VDD.n843 DVSS 0.082647f
C4159 VDD.n844 DVSS 0.082647f
C4160 VDD.n845 DVSS 0.01686f
C4161 VDD.n846 DVSS 0.02248f
C4162 VDD.n847 DVSS 0.026688f
C4163 VDD.n848 DVSS 0.055959f
C4164 VDD.t125 DVSS 0.038224f
C4165 VDD.t85 DVSS 0.028927f
C4166 VDD.n849 DVSS 0.079201f
C4167 VDD.n850 DVSS 0.013612f
C4168 VDD.n851 DVSS 0.210629f
C4169 VDD.n852 DVSS 0.068012f
C4170 VDD.n853 DVSS 0.068873f
C4171 VDD.n854 DVSS 0.02248f
C4172 VDD.n855 DVSS 0.02248f
C4173 VDD.n856 DVSS 0.02841f
C4174 VDD.n857 DVSS 0.02358f
C4175 VDD.t124 DVSS 0.028448f
C4176 VDD.n858 DVSS 0.049105f
C4177 VDD.n859 DVSS 1.32039f
C4178 VDD.n860 DVSS 0.055959f
C4179 VDD.n861 DVSS 0.037467f
C4180 VDD.n862 DVSS 0.02248f
C4181 VDD.n863 DVSS 0.082647f
C4182 VDD.n864 DVSS 0.041324f
C4183 VDD.n865 DVSS 0.129401f
C4184 VDD.n866 DVSS 0.170494f
C4185 VDD.n867 DVSS 0.088433f
C4186 VDD.n868 DVSS 0.041324f
C4187 VDD.n869 DVSS 0.062846f
C4188 VDD.n870 DVSS 0.02248f
C4189 VDD.n871 DVSS 0.01686f
C4190 VDD.n872 DVSS 0.082647f
C4191 VDD.n873 DVSS 0.082647f
C4192 VDD.n874 DVSS 0.01686f
C4193 VDD.n875 DVSS 0.02248f
C4194 VDD.n876 DVSS 0.026688f
C4195 VDD.n877 DVSS 0.055959f
C4196 VDD.t225 DVSS 0.038224f
C4197 VDD.t189 DVSS 0.028927f
C4198 VDD.n878 DVSS 0.079201f
C4199 VDD.n879 DVSS 0.013612f
C4200 VDD.n880 DVSS 0.210629f
C4201 VDD.n881 DVSS 0.068012f
C4202 VDD.n882 DVSS 0.068873f
C4203 VDD.n883 DVSS 0.02248f
C4204 VDD.n884 DVSS 0.02248f
C4205 VDD.n885 DVSS 0.02841f
C4206 VDD.n886 DVSS 0.02358f
C4207 VDD.t224 DVSS 0.028448f
C4208 VDD.n887 DVSS 0.049105f
C4209 VDD.n888 DVSS 1.32039f
C4210 VDD.n889 DVSS 0.055959f
C4211 VDD.n890 DVSS 0.037467f
C4212 VDD.n891 DVSS 0.02248f
C4213 VDD.n892 DVSS 0.082647f
C4214 VDD.n893 DVSS 0.041324f
C4215 VDD.n894 DVSS 0.129401f
C4216 VDD.n895 DVSS 0.170494f
C4217 VDD.n896 DVSS 0.088433f
C4218 VDD.n897 DVSS 0.041324f
C4219 VDD.n898 DVSS 0.062846f
C4220 VDD.n899 DVSS 0.02248f
C4221 VDD.n900 DVSS 0.01686f
C4222 VDD.n901 DVSS 0.082647f
C4223 VDD.n902 DVSS 0.082647f
C4224 VDD.n903 DVSS 0.01686f
C4225 VDD.n904 DVSS 0.02248f
C4226 VDD.n905 DVSS 0.026688f
C4227 VDD.n906 DVSS 0.055959f
C4228 VDD.t89 DVSS 0.038224f
C4229 VDD.t166 DVSS 0.028927f
C4230 VDD.n907 DVSS 0.079201f
C4231 VDD.n908 DVSS 0.013612f
C4232 VDD.n909 DVSS 0.210629f
C4233 VDD.n910 DVSS 0.068012f
C4234 VDD.n911 DVSS 0.068873f
C4235 VDD.n912 DVSS 0.02248f
C4236 VDD.n913 DVSS 0.02248f
C4237 VDD.n914 DVSS 0.02841f
C4238 VDD.n915 DVSS 0.02358f
C4239 VDD.t87 DVSS 0.028448f
C4240 VDD.n916 DVSS 0.049105f
C4241 VDD.n917 DVSS 1.32039f
C4242 VDD.n918 DVSS 0.055959f
C4243 VDD.n919 DVSS 0.037467f
C4244 VDD.n920 DVSS 0.02248f
C4245 VDD.n921 DVSS 0.082647f
C4246 VDD.n922 DVSS 0.041324f
C4247 VDD.n923 DVSS 0.129401f
C4248 VDD.n924 DVSS 0.170494f
C4249 VDD.n925 DVSS 0.088433f
C4250 VDD.n926 DVSS 0.041324f
C4251 VDD.n927 DVSS 0.062846f
C4252 VDD.n928 DVSS 0.02248f
C4253 VDD.n929 DVSS 0.01686f
C4254 VDD.n930 DVSS 0.082647f
C4255 VDD.n931 DVSS 0.082647f
C4256 VDD.n932 DVSS 0.01686f
C4257 VDD.n933 DVSS 0.02248f
C4258 VDD.n934 DVSS 0.026688f
C4259 VDD.n935 DVSS 0.055959f
C4260 VDD.t57 DVSS 0.038224f
C4261 VDD.t9 DVSS 0.028927f
C4262 VDD.n936 DVSS 0.079201f
C4263 VDD.n937 DVSS 0.013612f
C4264 VDD.n938 DVSS 0.210629f
C4265 VDD.n939 DVSS 0.068012f
C4266 VDD.n940 DVSS 0.068873f
C4267 VDD.n941 DVSS 0.02248f
C4268 VDD.n942 DVSS 0.02248f
C4269 VDD.n943 DVSS 0.02841f
C4270 VDD.n944 DVSS 0.02358f
C4271 VDD.t56 DVSS 0.028448f
C4272 VDD.n945 DVSS 0.049105f
C4273 VDD.n946 DVSS 1.32039f
C4274 VDD.n947 DVSS 0.055959f
C4275 VDD.n948 DVSS 0.037467f
C4276 VDD.n949 DVSS 0.02248f
C4277 VDD.n950 DVSS 0.082647f
C4278 VDD.n951 DVSS 0.041324f
C4279 VDD.n952 DVSS 0.129401f
C4280 VDD.n953 DVSS 0.170494f
C4281 VDD.n954 DVSS 0.088433f
C4282 VDD.n955 DVSS 0.041324f
C4283 VDD.n956 DVSS 0.062846f
C4284 VDD.n957 DVSS 0.02248f
C4285 VDD.n958 DVSS 0.01686f
C4286 VDD.n959 DVSS 0.082647f
C4287 VDD.n960 DVSS 0.082647f
C4288 VDD.n961 DVSS 0.01686f
C4289 VDD.n962 DVSS 0.02248f
C4290 VDD.n963 DVSS 0.026688f
C4291 VDD.n964 DVSS 0.055959f
C4292 VDD.t181 DVSS 0.038224f
C4293 VDD.t114 DVSS 0.028927f
C4294 VDD.n965 DVSS 0.079201f
C4295 VDD.n966 DVSS 0.013612f
C4296 VDD.n967 DVSS 0.210629f
C4297 VDD.n968 DVSS 0.068012f
C4298 VDD.n969 DVSS 0.068873f
C4299 VDD.n970 DVSS 0.02248f
C4300 VDD.n971 DVSS 0.02248f
C4301 VDD.n972 DVSS 0.02841f
C4302 VDD.n973 DVSS 0.02358f
C4303 VDD.t180 DVSS 0.028448f
C4304 VDD.n974 DVSS 0.049105f
C4305 VDD.n975 DVSS 1.32039f
C4306 VDD.n976 DVSS 0.055959f
C4307 VDD.n977 DVSS 0.037467f
C4308 VDD.n978 DVSS 0.02248f
C4309 VDD.n979 DVSS 0.082647f
C4310 VDD.n980 DVSS 0.041324f
C4311 VDD.n981 DVSS 0.129401f
C4312 VDD.n982 DVSS 0.170494f
C4313 VDD.n983 DVSS 0.088433f
C4314 VDD.n984 DVSS 0.041324f
C4315 VDD.n985 DVSS 0.062846f
C4316 VDD.n986 DVSS 0.02248f
C4317 VDD.n987 DVSS 0.01686f
C4318 VDD.n988 DVSS 0.082647f
C4319 VDD.n989 DVSS 0.082647f
C4320 VDD.n990 DVSS 0.01686f
C4321 VDD.n991 DVSS 0.02248f
C4322 VDD.n992 DVSS 0.026688f
C4323 VDD.n993 DVSS 0.055959f
C4324 VDD.t195 DVSS 0.038224f
C4325 VDD.t103 DVSS 0.028927f
C4326 VDD.n994 DVSS 0.079201f
C4327 VDD.n995 DVSS 0.013612f
C4328 VDD.n996 DVSS 0.210629f
C4329 VDD.n997 DVSS 0.068012f
C4330 VDD.n998 DVSS 0.068873f
C4331 VDD.n999 DVSS 0.02248f
C4332 VDD.n1000 DVSS 0.02248f
C4333 VDD.n1001 DVSS 0.02841f
C4334 VDD.n1002 DVSS 0.02358f
C4335 VDD.t197 DVSS 0.028448f
C4336 VDD.n1003 DVSS 0.049105f
C4337 VDD.n1004 DVSS 0.638554f
C4338 VDD.n1005 DVSS 2.17483f
C4339 VDD.n1006 DVSS 3.97069f
C4340 VDD.n1007 DVSS 29.399801f
C4341 a_1031_764.n0 DVSS 5.39149f
C4342 a_1031_764.n1 DVSS 1.18632f
C4343 a_1031_764.n2 DVSS 5.40279f
C4344 a_1031_764.t3 DVSS 0.194246f
C4345 a_1031_764.t7 DVSS 2.01847f
C4346 a_1031_764.n3 DVSS 0.484536f
C4347 a_1031_764.t4 DVSS 2.01847f
C4348 a_1031_764.n4 DVSS 0.016223f
C4349 a_1031_764.t6 DVSS 2.01847f
C4350 a_1031_764.n5 DVSS 0.017021f
C4351 a_1031_764.t5 DVSS 2.01847f
C4352 a_1031_764.n6 DVSS 1.56837f
C4353 a_1031_764.n7 DVSS 1.07807f
C4354 a_1031_764.t2 DVSS 10.7549f
C4355 a_1031_764.n8 DVSS 0.873302f
C4356 a_1031_764.t1 DVSS 1.68114f
C4357 a_1031_764.n9 DVSS 1.48738f
C4358 a_1031_764.n10 DVSS 0.396152f
C4359 a_1031_764.t0 DVSS 0.194246f
C4360 VSS.n0 DVSS 0.238708f
C4361 VSS.n1 DVSS 0.348086f
C4362 VSS.n2 DVSS 0.737969f
C4363 VSS.n3 DVSS 0.094511f
C4364 VSS.n4 DVSS 0.094511f
C4365 VSS.n5 DVSS 0.305052f
C4366 VSS.n6 DVSS 0.254689f
C4367 VSS.n7 DVSS 1.60661f
C4368 VSS.n8 DVSS 0.255534f
C4369 VSS.n9 DVSS 0.255534f
C4370 VSS.n10 DVSS 0.902438f
C4371 VSS.n11 DVSS 0.341966f
C4372 VSS.n12 DVSS 0.380541f
C4373 VSS.n13 DVSS 0.586221f
C4374 VSS.n14 DVSS 0.427512f
C4375 VSS.n15 DVSS 0.594373f
C4376 VSS.n16 DVSS 0.427512f
C4377 VSS.n17 DVSS 0.594373f
C4378 VSS.n18 DVSS 0.427512f
C4379 VSS.n19 DVSS 0.594373f
C4380 VSS.n20 DVSS 0.704567f
C4381 VSS.n21 DVSS 0.697161f
C4382 VSS.n22 DVSS 0.597705f
C4383 VSS.n23 DVSS 0.135668f
C4384 VSS.n24 DVSS 0.317221f
C4385 VSS.n25 DVSS 0.285633f
C4386 VSS.n26 DVSS 0.285633f
C4387 VSS.t245 DVSS 2.62345f
C4388 VSS.n27 DVSS 0.282707f
C4389 VSS.n28 DVSS 0.282707f
C4390 VSS.n29 DVSS 0.569431f
C4391 VSS.n30 DVSS 0.285633f
C4392 VSS.n31 DVSS 0.285633f
C4393 VSS.n32 DVSS 0.518818f
C4394 VSS.n33 DVSS 0.862405f
C4395 VSS.n34 DVSS 0.255534f
C4396 VSS.n35 DVSS 0.025874f
C4397 VSS.n36 DVSS 2.37941f
C4398 VSS.n37 DVSS 3.17255f
C4399 VSS.n38 DVSS 0.36621f
C4400 VSS.n39 DVSS 0.482775f
C4401 VSS.n40 DVSS 0.244293f
C4402 VSS.n41 DVSS 0.277011f
C4403 VSS.n42 DVSS 0.277011f
C4404 VSS.n43 DVSS 0.277011f
C4405 VSS.n44 DVSS 0.505013f
C4406 VSS.n45 DVSS 0.128365f
C4407 VSS.n46 DVSS 0.206917f
C4408 VSS.n47 DVSS 0.206917f
C4409 VSS.t58 DVSS 2.62345f
C4410 VSS.n48 DVSS 0.206767f
C4411 VSS.n49 DVSS 0.206767f
C4412 VSS.n50 DVSS 1.66762f
C4413 VSS.n51 DVSS 0.206917f
C4414 VSS.n52 DVSS 0.206917f
C4415 VSS.n53 DVSS 0.421535f
C4416 VSS.n54 DVSS 0.593348f
C4417 VSS.n55 DVSS 0.210893f
C4418 VSS.n56 DVSS 0.212563f
C4419 VSS.n57 DVSS 0.053507f
C4420 VSS.t75 DVSS 3.7013f
C4421 VSS.t167 DVSS 2.11503f
C4422 VSS.n58 DVSS 0.66183f
C4423 VSS.n59 DVSS 0.212563f
C4424 VSS.n60 DVSS 2.06501f
C4425 VSS.n61 DVSS 0.014658f
C4426 VSS.n62 DVSS 0.267615f
C4427 VSS.n63 DVSS 0.286553f
C4428 VSS.n64 DVSS 0.286553f
C4429 VSS.n65 DVSS 0.286553f
C4430 VSS.n66 DVSS 0.552922f
C4431 VSS.n67 DVSS 0.054985f
C4432 VSS.n68 DVSS 0.168383f
C4433 VSS.n69 DVSS 0.168383f
C4434 VSS.t99 DVSS 2.62345f
C4435 VSS.n70 DVSS 0.170661f
C4436 VSS.n71 DVSS 0.170661f
C4437 VSS.n72 DVSS 2.62345f
C4438 VSS.n73 DVSS 0.168383f
C4439 VSS.n74 DVSS 0.168383f
C4440 VSS.n75 DVSS 0.277508f
C4441 VSS.n76 DVSS 0.584036f
C4442 VSS.n77 DVSS 0.188923f
C4443 VSS.n78 DVSS 0.191148f
C4444 VSS.n79 DVSS 0.08234f
C4445 VSS.t192 DVSS 3.82332f
C4446 VSS.n80 DVSS 1.52526f
C4447 VSS.n81 DVSS 0.191148f
C4448 VSS.n82 DVSS 0.191148f
C4449 VSS.n83 DVSS 0.223152f
C4450 VSS.n84 DVSS 0.180466f
C4451 VSS.n85 DVSS 0.180466f
C4452 VSS.n86 DVSS 3.19288f
C4453 VSS.n87 DVSS 0.177913f
C4454 VSS.t119 DVSS 2.09469f
C4455 VSS.n88 DVSS 0.178319f
C4456 VSS.n89 DVSS 0.201105f
C4457 VSS.n90 DVSS 0.31291f
C4458 VSS.n91 DVSS 0.456818f
C4459 VSS.n92 DVSS 0.398407f
C4460 VSS.n93 DVSS 0.246725f
C4461 VSS.n94 DVSS 0.324725f
C4462 VSS.n95 DVSS 0.210354f
C4463 VSS.t182 DVSS 0.345726f
C4464 VSS.n96 DVSS 5.14522f
C4465 VSS.n97 DVSS 0.210354f
C4466 VSS.n98 DVSS 0.053941f
C4467 VSS.n99 DVSS 0.212638f
C4468 VSS.n100 DVSS 0.737969f
C4469 VSS.n101 DVSS 0.324725f
C4470 VSS.n102 DVSS 0.335946f
C4471 VSS.n103 DVSS 5.75532f
C4472 VSS.n104 DVSS 0.284716f
C4473 VSS.n105 DVSS 0.074079f
C4474 VSS.n106 DVSS 0.376118f
C4475 VSS.n107 DVSS 0.376118f
C4476 VSS.t9 DVSS 4.51478f
C4477 VSS.t47 DVSS 2.15432f
C4478 VSS.n108 DVSS 0.949994f
C4479 VSS.t70 DVSS 0.506969f
C4480 VSS.n109 DVSS 1.6765f
C4481 VSS.n110 DVSS 4.9285f
C4482 VSS.n111 DVSS 5.71627f
C4483 VSS.t219 DVSS 0.412654f
C4484 VSS.n112 DVSS 1.2573f
C4485 VSS.n113 DVSS 0.981055f
C4486 VSS.n114 DVSS 0.080615f
C4487 VSS.n115 DVSS 0.523872f
C4488 VSS.n116 DVSS 0.201105f
C4489 VSS.n117 DVSS 0.31291f
C4490 VSS.n118 DVSS 1.05752f
C4491 VSS.t72 DVSS 1.56594f
C4492 VSS.n119 DVSS 0.200927f
C4493 VSS.n120 DVSS 0.132568f
C4494 VSS.n121 DVSS 0.053941f
C4495 VSS.n122 DVSS 0.398407f
C4496 VSS.n123 DVSS 0.184271f
C4497 VSS.n124 DVSS 0.184271f
C4498 VSS.t48 DVSS 3.96568f
C4499 VSS.n125 DVSS 4.57579f
C4500 VSS.t28 DVSS 1.46425f
C4501 VSS.t196 DVSS 1.68796f
C4502 VSS.t171 DVSS 3.19288f
C4503 VSS.n126 DVSS 0.094511f
C4504 VSS.n127 DVSS 0.096637f
C4505 VSS.n128 DVSS 0.153316f
C4506 VSS.n129 DVSS 1.932f
C4507 VSS.t208 DVSS 4.14871f
C4508 VSS.n130 DVSS 0.376118f
C4509 VSS.n131 DVSS 0.376118f
C4510 VSS.n132 DVSS 0.763628f
C4511 VSS.n133 DVSS 0.055762f
C4512 VSS.n134 DVSS 0.206313f
C4513 VSS.n135 DVSS 0.210354f
C4514 VSS.n136 DVSS 0.324725f
C4515 VSS.t108 DVSS 3.66063f
C4516 VSS.t197 DVSS 4.2504f
C4517 VSS.t3 DVSS 3.72164f
C4518 VSS.n137 DVSS 0.210354f
C4519 VSS.t34 DVSS 4.12838f
C4520 VSS.t55 DVSS 2.86749f
C4521 VSS.t31 DVSS 4.02669f
C4522 VSS.n138 DVSS 3.11153f
C4523 VSS.n139 DVSS 0.335946f
C4524 VSS.n140 DVSS 0.212638f
C4525 VSS.n141 DVSS 0.154979f
C4526 VSS.n142 DVSS 0.246725f
C4527 VSS.n143 DVSS 0.949994f
C4528 VSS.n144 DVSS 0.456818f
C4529 VSS.n145 DVSS 0.31291f
C4530 VSS.n146 DVSS 0.201105f
C4531 VSS.t200 DVSS 2.60311f
C4532 VSS.t89 DVSS 3.76231f
C4533 VSS.n147 DVSS 0.200927f
C4534 VSS.n148 DVSS 1.6765f
C4535 VSS.t50 DVSS 0.412654f
C4536 VSS.n149 DVSS 1.2573f
C4537 VSS.n150 DVSS 0.096637f
C4538 VSS.n151 DVSS 0.616198f
C4539 VSS.n152 DVSS 0.31291f
C4540 VSS.t153 DVSS 2.7048f
C4541 VSS.n153 DVSS 0.317213f
C4542 VSS.n154 DVSS 2.3184f
C4543 VSS.n155 DVSS 2.5421f
C4544 VSS.t88 DVSS 2.44042f
C4545 VSS.t151 DVSS 2.62345f
C4546 VSS.n156 DVSS 2.35907f
C4547 VSS.n157 DVSS 2.25739f
C4548 VSS.n158 DVSS 0.398407f
C4549 VSS.n159 DVSS 0.246725f
C4550 VSS.n160 DVSS 0.391577f
C4551 VSS.n161 DVSS 0.324725f
C4552 VSS.n162 DVSS 0.210354f
C4553 VSS.t159 DVSS 0.711789f
C4554 VSS.t32 DVSS 4.81983f
C4555 VSS.n163 DVSS 0.210354f
C4556 VSS.n164 DVSS 0.053941f
C4557 VSS.n165 DVSS 0.212638f
C4558 VSS.n166 DVSS 0.737969f
C4559 VSS.n167 DVSS 0.324725f
C4560 VSS.n168 DVSS 3.7013f
C4561 VSS.n169 DVSS 4.18939f
C4562 VSS.n170 DVSS 0.122364f
C4563 VSS.n171 DVSS 0.376118f
C4564 VSS.n172 DVSS 0.376118f
C4565 VSS.t71 DVSS 3.27423f
C4566 VSS.n173 DVSS 0.206767f
C4567 VSS.n174 DVSS 0.206767f
C4568 VSS.n175 DVSS 0.752463f
C4569 VSS.n176 DVSS 0.206767f
C4570 VSS.n177 DVSS 0.206917f
C4571 VSS.n178 DVSS 0.206917f
C4572 VSS.n179 DVSS 0.421535f
C4573 VSS.n180 DVSS 0.593348f
C4574 VSS.n181 DVSS 0.210893f
C4575 VSS.n182 DVSS 0.212563f
C4576 VSS.n183 DVSS 0.032718f
C4577 VSS.n184 DVSS 3.23356f
C4578 VSS.n185 DVSS 0.210893f
C4579 VSS.n186 DVSS 0.206917f
C4580 VSS.n187 DVSS 2.74547f
C4581 VSS.n188 DVSS 0.178407f
C4582 VSS.n189 DVSS 0.31291f
C4583 VSS.n190 DVSS 0.201105f
C4584 VSS.n191 DVSS 0.997699f
C4585 VSS.n192 DVSS 0.116656f
C4586 VSS.t74 DVSS 0.412654f
C4587 VSS.n193 DVSS 1.2573f
C4588 VSS.t207 DVSS 0.412654f
C4589 VSS.n194 DVSS 1.02936f
C4590 VSS.n195 DVSS 0.294032f
C4591 VSS.n196 DVSS 4.9285f
C4592 VSS.n197 DVSS 5.71627f
C4593 VSS.n198 DVSS 5.87937f
C4594 VSS.n199 DVSS 6.77815f
C4595 VSS.n200 DVSS 0.165495f
C4596 VSS.n201 DVSS 0.210152f
C4597 VSS.n202 DVSS 0.10449f
C4598 VSS.n203 DVSS 0.145623f
C4599 VSS.t163 DVSS 3.84366f
C4600 VSS.n204 DVSS 0.093231f
C4601 VSS.t115 DVSS 3.55895f
C4602 VSS.n205 DVSS 0.093231f
C4603 VSS.n206 DVSS 0.10449f
C4604 VSS.n207 DVSS 0.145623f
C4605 VSS.n208 DVSS 0.036109f
C4606 VSS.n209 DVSS 0.206373f
C4607 VSS.n210 DVSS 0.082794f
C4608 VSS.n211 DVSS 0.042179f
C4609 VSS.n212 DVSS 0.348559f
C4610 VSS.n213 DVSS 0.197943f
C4611 VSS.n214 DVSS 0.197943f
C4612 VSS.n215 DVSS 0.197943f
C4613 VSS.n216 DVSS 0.197943f
C4614 VSS.n217 DVSS 0.156375f
C4615 VSS.n218 DVSS 0.180466f
C4616 VSS.n219 DVSS 0.180466f
C4617 VSS.n220 DVSS 1.80998f
C4618 VSS.n221 DVSS 0.180466f
C4619 VSS.n222 DVSS 0.180466f
C4620 VSS.n223 DVSS 0.082547f
C4621 VSS.n224 DVSS 0.185526f
C4622 VSS.n225 DVSS 0.197943f
C4623 VSS.n226 DVSS 0.197943f
C4624 VSS.n227 DVSS 0.286553f
C4625 VSS.n228 DVSS 0.552922f
C4626 VSS.n229 DVSS 0.03485f
C4627 VSS.n230 DVSS 0.032827f
C4628 VSS.n231 DVSS 0.343189f
C4629 VSS.n232 DVSS 0.10449f
C4630 VSS.n233 DVSS 5.32825f
C4631 VSS.n234 DVSS 0.124219f
C4632 VSS.n235 DVSS 5.38926f
C4633 VSS.n236 DVSS 0.210354f
C4634 VSS.n237 DVSS 0.210354f
C4635 VSS.n238 DVSS 0.246725f
C4636 VSS.n239 DVSS 0.055762f
C4637 VSS.n240 DVSS 0.210362f
C4638 VSS.n241 DVSS 0.184271f
C4639 VSS.n242 DVSS 0.354664f
C4640 VSS.n243 DVSS 0.280181f
C4641 VSS.n244 DVSS 56.5667f
C4642 VSS.n245 DVSS 0.094511f
C4643 VSS.n246 DVSS 0.094511f
C4644 VSS.n247 DVSS 0.949994f
C4645 VSS.t136 DVSS 0.506969f
C4646 VSS.t135 DVSS 2.35907f
C4647 VSS.t120 DVSS 1.89133f
C4648 VSS.t127 DVSS 3.4776f
C4649 VSS.t123 DVSS 2.27587f
C4650 VSS.t226 DVSS 1.76728f
C4651 VSS.n248 DVSS 4.75882f
C4652 VSS.n249 DVSS 0.369019f
C4653 VSS.n250 DVSS 1.54772f
C4654 VSS.n251 DVSS 1.67792f
C4655 VSS.n252 DVSS 0.018952f
C4656 VSS.n253 DVSS 0.129233f
C4657 VSS.n254 DVSS 0.671674f
C4658 VSS.n255 DVSS 0.277011f
C4659 VSS.n256 DVSS 0.277011f
C4660 VSS.n257 DVSS 0.277011f
C4661 VSS.n258 DVSS 0.277011f
C4662 VSS.n259 DVSS 0.224526f
C4663 VSS.n260 DVSS 0.046972f
C4664 VSS.n261 DVSS 0.380541f
C4665 VSS.n262 DVSS 0.014658f
C4666 VSS.n263 DVSS 0.267615f
C4667 VSS.n264 DVSS 0.286553f
C4668 VSS.n265 DVSS 0.286553f
C4669 VSS.n266 DVSS 0.054985f
C4670 VSS.n267 DVSS 0.168383f
C4671 VSS.n268 DVSS 0.168383f
C4672 VSS.t241 DVSS 2.35907f
C4673 VSS.n269 DVSS 0.170661f
C4674 VSS.n270 DVSS 0.170661f
C4675 VSS.n271 DVSS 2.44042f
C4676 VSS.n272 DVSS 0.168383f
C4677 VSS.n273 DVSS 0.168383f
C4678 VSS.n274 DVSS 0.277508f
C4679 VSS.n275 DVSS 0.584036f
C4680 VSS.n276 DVSS 0.188923f
C4681 VSS.n277 DVSS 0.191148f
C4682 VSS.n278 DVSS 0.08234f
C4683 VSS.t41 DVSS 3.84366f
C4684 VSS.n279 DVSS 1.50493f
C4685 VSS.n280 DVSS 0.191148f
C4686 VSS.n281 DVSS 0.191148f
C4687 VSS.n282 DVSS 0.223152f
C4688 VSS.n283 DVSS 0.180466f
C4689 VSS.n284 DVSS 0.10606f
C4690 VSS.n285 DVSS 0.286553f
C4691 VSS.n286 DVSS 0.10606f
C4692 VSS.n287 DVSS 0.286553f
C4693 VSS.n288 DVSS 0.10606f
C4694 VSS.n289 DVSS 0.286553f
C4695 VSS.n290 DVSS 0.10606f
C4696 VSS.n291 DVSS 0.286553f
C4697 VSS.n292 DVSS 0.221965f
C4698 VSS.n293 DVSS 0.489521f
C4699 VSS.n294 DVSS 0.112492f
C4700 VSS.n295 DVSS 0.114447f
C4701 VSS.n296 DVSS 0.13796f
C4702 VSS.n297 DVSS 0.13796f
C4703 VSS.n298 DVSS 0.13796f
C4704 VSS.n299 DVSS 0.13796f
C4705 VSS.n300 DVSS 0.273916f
C4706 VSS.n301 DVSS 0.11972f
C4707 VSS.n302 DVSS 0.343918f
C4708 VSS.n303 DVSS 0.02564f
C4709 VSS.n304 DVSS 0.228351f
C4710 VSS.n305 DVSS 0.331014f
C4711 VSS.n306 DVSS 0.197943f
C4712 VSS.n307 DVSS 0.197943f
C4713 VSS.n308 DVSS 0.197943f
C4714 VSS.n309 DVSS 0.197943f
C4715 VSS.n310 DVSS 0.156375f
C4716 VSS.n311 DVSS 0.177913f
C4717 VSS.n312 DVSS 0.053984f
C4718 VSS.n313 DVSS 0.177913f
C4719 VSS.n314 DVSS 0.180466f
C4720 VSS.n315 DVSS 1.66762f
C4721 VSS.n316 DVSS 0.177913f
C4722 VSS.n317 DVSS 0.10449f
C4723 VSS.n318 DVSS 0.093231f
C4724 VSS.n319 DVSS 0.093231f
C4725 VSS.n320 DVSS 0.184271f
C4726 VSS.n321 DVSS 0.324725f
C4727 VSS.n322 DVSS 0.391577f
C4728 VSS.n323 DVSS 0.178319f
C4729 VSS.n324 DVSS 0.200927f
C4730 VSS.n325 DVSS 0.253124f
C4731 VSS.n326 DVSS 0.370974f
C4732 VSS.n327 DVSS 0.188923f
C4733 VSS.n328 DVSS 4.88084f
C4734 VSS.n329 DVSS 0.317213f
C4735 VSS.n330 DVSS 3.07086f
C4736 VSS.t154 DVSS 0.732126f
C4737 VSS.n331 DVSS 0.630442f
C4738 VSS.n332 DVSS 0.096637f
C4739 VSS.n333 DVSS 0.132568f
C4740 VSS.n334 DVSS 0.053941f
C4741 VSS.n335 DVSS 0.616198f
C4742 VSS.n336 DVSS 0.256757f
C4743 VSS.t155 DVSS 0.325389f
C4744 VSS.t133 DVSS 2.23705f
C4745 VSS.n337 DVSS 0.178319f
C4746 VSS.n338 DVSS 0.31291f
C4747 VSS.n339 DVSS 0.398407f
C4748 VSS.n340 DVSS 0.532664f
C4749 VSS.n341 DVSS 0.154979f
C4750 VSS.n342 DVSS 0.184271f
C4751 VSS.t122 DVSS 3.72164f
C4752 VSS.n343 DVSS 0.093231f
C4753 VSS.n344 DVSS 0.145623f
C4754 VSS.n345 DVSS 0.031491f
C4755 VSS.n346 DVSS 0.057447f
C4756 VSS.n347 DVSS 0.20043f
C4757 VSS.n348 DVSS 0.263852f
C4758 VSS.n349 DVSS 0.13796f
C4759 VSS.n350 DVSS 0.13796f
C4760 VSS.n351 DVSS 0.13796f
C4761 VSS.n352 DVSS 0.13796f
C4762 VSS.n353 DVSS 0.223503f
C4763 VSS.n354 DVSS 0.200056f
C4764 VSS.n355 DVSS 0.211575f
C4765 VSS.n356 DVSS 0.211575f
C4766 VSS.n357 DVSS 0.211575f
C4767 VSS.n358 DVSS 0.421535f
C4768 VSS.n359 DVSS 0.341419f
C4769 VSS.n360 DVSS 0.128365f
C4770 VSS.n361 DVSS 0.12758f
C4771 VSS.n362 DVSS 1.14874f
C4772 VSS.n363 DVSS 0.285633f
C4773 VSS.n364 DVSS 0.518818f
C4774 VSS.n365 DVSS 0.206917f
C4775 VSS.n366 DVSS 0.136864f
C4776 VSS.n367 DVSS 0.862405f
C4777 VSS.n368 DVSS 0.254689f
C4778 VSS.n369 DVSS 0.255534f
C4779 VSS.n370 DVSS 0.025874f
C4780 VSS.t124 DVSS 1.85065f
C4781 VSS.n371 DVSS 0.335946f
C4782 VSS.n372 DVSS 2.37941f
C4783 VSS.n373 DVSS 0.255534f
C4784 VSS.n374 DVSS 0.254689f
C4785 VSS.n375 DVSS 0.311212f
C4786 VSS.n376 DVSS 0.704567f
C4787 VSS.n377 DVSS 0.659377f
C4788 VSS.n378 DVSS 0.282707f
C4789 VSS.n379 DVSS 0.285633f
C4790 VSS.n380 DVSS 0.367012f
C4791 VSS.n381 DVSS 0.129985f
C4792 VSS.n382 DVSS 0.649633f
C4793 VSS.n383 DVSS 0.571907f
C4794 VSS.n384 DVSS 0.427512f
C4795 VSS.n385 DVSS 0.54257f
C4796 VSS.n386 DVSS 0.427512f
C4797 VSS.n387 DVSS 0.54257f
C4798 VSS.n388 DVSS 0.427512f
C4799 VSS.n389 DVSS 0.54257f
C4800 VSS.n390 DVSS 0.427512f
C4801 VSS.n391 DVSS 0.54257f
C4802 VSS.n392 DVSS 0.36621f
C4803 VSS.n393 DVSS 0.526211f
C4804 VSS.n394 DVSS 0.341966f
C4805 VSS.n395 DVSS 0.401638f
C4806 VSS.n396 DVSS 0.016768f
C4807 VSS.n397 DVSS 0.54257f
C4808 VSS.n398 DVSS 0.427512f
C4809 VSS.n399 DVSS 0.54257f
C4810 VSS.n400 DVSS 0.427512f
C4811 VSS.n401 DVSS 0.54257f
C4812 VSS.n402 DVSS 0.427512f
C4813 VSS.n403 DVSS 0.54257f
C4814 VSS.n404 DVSS 0.704567f
C4815 VSS.n405 DVSS 0.576924f
C4816 VSS.n406 DVSS 0.602989f
C4817 VSS.n407 DVSS 0.341792f
C4818 VSS.t172 DVSS 5.06387f
C4819 VSS.n408 DVSS 0.341792f
C4820 VSS.n409 DVSS 0.341792f
C4821 VSS.n410 DVSS 0.536899f
C4822 VSS.n411 DVSS 0.110398f
C4823 VSS.n412 DVSS 0.951024f
C4824 VSS.n413 DVSS 0.971718f
C4825 VSS.n414 DVSS 0.971718f
C4826 VSS.n415 DVSS 0.427512f
C4827 VSS.n416 DVSS 0.427512f
C4828 VSS.n417 DVSS 0.427512f
C4829 VSS.n418 DVSS 0.971718f
C4830 VSS.n419 DVSS 1.28393f
C4831 VSS.n420 DVSS 0.061871f
C4832 VSS.n421 DVSS 0.597705f
C4833 VSS.n422 DVSS 0.409292f
C4834 VSS.n423 DVSS 0.999855f
C4835 VSS.n424 DVSS 0.518818f
C4836 VSS.n425 DVSS 0.135668f
C4837 VSS.n426 DVSS 0.409292f
C4838 VSS.t103 DVSS 3.29457f
C4839 VSS.n427 DVSS 0.370974f
C4840 VSS.n428 DVSS 0.253124f
C4841 VSS.n429 DVSS 0.178407f
C4842 VSS.t105 DVSS 3.19039f
C4843 VSS.t18 DVSS 3.33524f
C4844 VSS.n430 DVSS 3.4776f
C4845 VSS.n431 DVSS 0.31291f
C4846 VSS.n432 DVSS 0.178319f
C4847 VSS.t218 DVSS 3.96568f
C4848 VSS.t223 DVSS 2.74547f
C4849 VSS.t138 DVSS 3.39625f
C4850 VSS.n433 DVSS 0.317213f
C4851 VSS.n434 DVSS 3.33524f
C4852 VSS.n435 DVSS 1.85065f
C4853 VSS.t54 DVSS 1.42358f
C4854 VSS.t183 DVSS 2.62345f
C4855 VSS.n436 DVSS 0.404475f
C4856 VSS.n437 DVSS 0.404475f
C4857 VSS.n438 DVSS 0.659421f
C4858 VSS.n439 DVSS 0.213335f
C4859 VSS.n440 DVSS 0.025193f
C4860 VSS.n441 DVSS 0.210152f
C4861 VSS.n442 DVSS 0.10449f
C4862 VSS.n443 DVSS 0.093231f
C4863 VSS.n444 DVSS 0.093231f
C4864 VSS.n445 DVSS 0.093231f
C4865 VSS.n446 DVSS 0.079713f
C4866 VSS.n447 DVSS 0.361477f
C4867 VSS.n448 DVSS 0.51729f
C4868 VSS.n449 DVSS 0.193204f
C4869 VSS.n450 DVSS 0.348559f
C4870 VSS.n451 DVSS 0.197943f
C4871 VSS.n452 DVSS 0.197943f
C4872 VSS.n453 DVSS 0.197943f
C4873 VSS.n454 DVSS 0.197943f
C4874 VSS.n455 DVSS 0.156375f
C4875 VSS.n456 DVSS 0.099037f
C4876 VSS.n457 DVSS 0.180466f
C4877 VSS.n458 DVSS 0.177913f
C4878 VSS.n459 DVSS 0.036109f
C4879 VSS.t173 DVSS 3.7013f
C4880 VSS.n460 DVSS 0.180466f
C4881 VSS.n461 DVSS 0.177913f
C4882 VSS.n462 DVSS 0.177913f
C4883 VSS.n463 DVSS 0.228351f
C4884 VSS.n464 DVSS 0.331014f
C4885 VSS.n465 DVSS 0.197943f
C4886 VSS.n466 DVSS 0.197943f
C4887 VSS.n467 DVSS 0.197943f
C4888 VSS.n468 DVSS 0.114447f
C4889 VSS.n469 DVSS 0.13796f
C4890 VSS.n470 DVSS 0.13796f
C4891 VSS.n471 DVSS 0.13796f
C4892 VSS.n472 DVSS 0.13796f
C4893 VSS.n473 DVSS 0.273916f
C4894 VSS.n474 DVSS 0.02564f
C4895 VSS.n475 DVSS 0.11972f
C4896 VSS.n476 DVSS 0.343918f
C4897 VSS.n477 DVSS 0.489521f
C4898 VSS.n478 DVSS 0.286553f
C4899 VSS.n479 DVSS 0.286553f
C4900 VSS.n480 DVSS 0.286553f
C4901 VSS.n481 DVSS 0.286553f
C4902 VSS.n482 DVSS 0.197943f
C4903 VSS.n483 DVSS 0.177913f
C4904 VSS.n484 DVSS 0.089876f
C4905 VSS.n485 DVSS 0.10606f
C4906 VSS.n486 DVSS 0.10606f
C4907 VSS.n487 DVSS 0.10606f
C4908 VSS.n488 DVSS 0.206373f
C4909 VSS.n489 DVSS 0.03485f
C4910 VSS.n490 DVSS 0.039888f
C4911 VSS.n491 DVSS 0.032827f
C4912 VSS.n492 DVSS 0.343189f
C4913 VSS.n493 DVSS 0.10449f
C4914 VSS.n494 DVSS 0.10449f
C4915 VSS.n495 DVSS 2.07436f
C4916 VSS.n496 DVSS 0.10449f
C4917 VSS.n497 DVSS 0.03485f
C4918 VSS.n498 DVSS 0.03464f
C4919 VSS.n499 DVSS 0.024186f
C4920 VSS.n500 DVSS 0.011288f
C4921 VSS.n501 DVSS 0.19695f
C4922 VSS.n502 DVSS 0.206373f
C4923 VSS.n503 DVSS 0.552922f
C4924 VSS.n504 DVSS 0.10606f
C4925 VSS.n505 DVSS 0.286553f
C4926 VSS.n506 DVSS 0.10606f
C4927 VSS.n507 DVSS 0.286553f
C4928 VSS.n508 DVSS 0.10606f
C4929 VSS.n509 DVSS 0.286553f
C4930 VSS.n510 DVSS 0.267615f
C4931 VSS.n511 DVSS 0.057447f
C4932 VSS.n512 DVSS 0.20043f
C4933 VSS.n513 DVSS 0.263852f
C4934 VSS.n514 DVSS 0.13796f
C4935 VSS.n515 DVSS 0.13796f
C4936 VSS.n516 DVSS 0.13796f
C4937 VSS.n517 DVSS 0.13796f
C4938 VSS.n518 DVSS 0.13796f
C4939 VSS.n519 DVSS 0.13796f
C4940 VSS.n520 DVSS 0.13796f
C4941 VSS.n521 DVSS 0.130937f
C4942 VSS.n522 DVSS 0.023971f
C4943 VSS.n523 DVSS 0.951024f
C4944 VSS.n524 DVSS 0.971718f
C4945 VSS.n525 DVSS 0.971718f
C4946 VSS.n526 DVSS 0.971718f
C4947 VSS.n527 DVSS 0.697161f
C4948 VSS.n528 DVSS 0.616976f
C4949 VSS.n529 DVSS 0.341966f
C4950 VSS.n530 DVSS 0.341966f
C4951 VSS.n531 DVSS 2.37941f
C4952 VSS.n532 DVSS 0.341792f
C4953 VSS.t188 DVSS 2.37941f
C4954 VSS.n533 DVSS 0.341792f
C4955 VSS.n534 DVSS 0.341966f
C4956 VSS.n535 DVSS 2.03551f
C4957 VSS.n536 DVSS 4.26694f
C4958 VSS.n537 DVSS 4.24175f
C4959 VSS.n538 DVSS 4.26854f
C4960 VSS.n539 DVSS 0.512401f
C4961 VSS.n540 DVSS 0.861497f
C4962 VSS.t199 DVSS 6.48999f
C4963 VSS.n541 DVSS 0.160742f
C4964 VSS.t235 DVSS 5.57687f
C4965 VSS.n542 DVSS 0.379528f
C4966 VSS.t215 DVSS 4.14251f
C4967 VSS.t169 DVSS 5.57687f
C4968 VSS.t237 DVSS 4.14251f
C4969 VSS.n543 DVSS 2.76168f
C4970 VSS.n544 DVSS 0.379528f
C4971 VSS.n545 DVSS 0.68552f
C4972 VSS.n546 DVSS 0.636296f
C4973 VSS.t216 DVSS 0.122081f
C4974 VSS.t238 DVSS 0.122081f
C4975 VSS.n547 DVSS 0.3828f
C4976 VSS.n548 DVSS 6.70272f
C4977 VSS.n549 DVSS 3.57924f
C4978 VSS.n550 DVSS 0.598752f
C4979 VSS.n551 DVSS 0.375413f
C4980 VSS.n552 DVSS 0.811402f
C4981 VSS.n553 DVSS 0.356133f
C4982 VSS.n554 DVSS 0.82035f
C4983 VSS.n555 DVSS 0.375413f
C4984 VSS.n556 DVSS 13.4692f
C4985 VSS.n557 DVSS 0.861497f
C4986 VSS.n558 DVSS 0.512401f
C4987 VSS.n559 DVSS 4.26654f
C4988 VSS.n560 DVSS 4.28903f
C4989 VSS.n561 DVSS 4.3872f
C4990 VSS.n562 DVSS 14.5023f
C4991 VSS.n563 DVSS 7.60646f
C4992 VSS.n564 DVSS 6.66772f
C4993 VSS.n565 DVSS 3.58831f
C4994 VSS.n566 DVSS 4.38665f
C4995 VSS.n567 DVSS 4.28903f
C4996 VSS.n568 DVSS 4.28957f
C4997 VSS.n569 DVSS 4.26708f
C4998 VSS.n570 DVSS 0.044987f
C4999 VSS.n571 DVSS 4.3907f
C5000 VSS.n572 DVSS 4.38827f
C5001 VSS.n573 DVSS 0.885933f
C5002 VSS.n574 DVSS 0.512401f
C5003 VSS.t102 DVSS 5.47349f
C5004 VSS.t51 DVSS 7.30124f
C5005 VSS.t29 DVSS 7.30124f
C5006 VSS.t42 DVSS 7.30124f
C5007 VSS.t57 DVSS 7.30124f
C5008 VSS.t112 DVSS 7.29794f
C5009 VSS.t184 DVSS 7.30051f
C5010 VSS.t30 DVSS 7.30124f
C5011 VSS.t116 DVSS 7.30124f
C5012 VSS.t60 DVSS 7.30124f
C5013 VSS.t77 DVSS 7.30124f
C5014 VSS.t39 DVSS 7.30124f
C5015 VSS.t79 DVSS 7.30124f
C5016 VSS.t141 DVSS 7.30124f
C5017 VSS.t174 DVSS 7.30124f
C5018 VSS.t91 DVSS 7.30124f
C5019 VSS.t0 DVSS 7.30124f
C5020 VSS.t160 DVSS 7.30124f
C5021 VSS.t118 DVSS 7.30038f
C5022 VSS.t6 DVSS 7.29808f
C5023 VSS.t104 DVSS 7.30124f
C5024 VSS.t4 DVSS 7.30124f
C5025 VSS.t145 DVSS 7.30124f
C5026 VSS.t126 DVSS 7.30124f
C5027 VSS.t13 DVSS 7.30124f
C5028 VSS.t43 DVSS 7.30124f
C5029 VSS.t143 DVSS 7.30124f
C5030 VSS.t8 DVSS 7.30124f
C5031 VSS.t150 DVSS 7.30124f
C5032 VSS.t157 DVSS 7.30124f
C5033 VSS.t40 DVSS 7.30124f
C5034 VSS.t27 DVSS 5.47593f
C5035 VSS.n575 DVSS 0.512401f
C5036 VSS.n576 DVSS 1.38139f
C5037 VSS.n577 DVSS 4.39128f
C5038 VSS.n578 DVSS 4.36569f
C5039 VSS.n579 DVSS 4.26906f
C5040 VSS.n580 DVSS 4.393f
C5041 VSS.n581 DVSS 4.2893f
C5042 VSS.n582 DVSS 4.2893f
C5043 VSS.n583 DVSS 4.38649f
C5044 VSS.n584 DVSS 4.28821f
C5045 VSS.n585 DVSS 4.26809f
C5046 VSS.n586 DVSS 0.044714f
C5047 VSS.n587 DVSS 4.28821f
C5048 VSS.n588 DVSS 4.26362f
C5049 VSS.n589 DVSS 4.26456f
C5050 VSS.n590 DVSS 0.044987f
C5051 VSS.n591 DVSS 0.160742f
C5052 VSS.t81 DVSS 3.35558f
C5053 VSS.t179 DVSS 5.14522f
C5054 VSS.n592 DVSS 0.376118f
C5055 VSS.n593 DVSS 0.369019f
C5056 VSS.n594 DVSS 0.369019f
C5057 VSS.n595 DVSS 0.20444f
C5058 VSS.n596 DVSS 0.080615f
C5059 VSS.t110 DVSS 0.506969f
C5060 VSS.n597 DVSS 1.56295f
C5061 VSS.n598 DVSS 0.178319f
C5062 VSS.n599 DVSS 0.200927f
C5063 VSS.n600 DVSS 0.256513f
C5064 VSS.n601 DVSS 1.94064f
C5065 VSS.t189 DVSS 0.412654f
C5066 VSS.n602 DVSS 1.2573f
C5067 VSS.n603 DVSS 0.096637f
C5068 VSS.n604 DVSS 0.616198f
C5069 VSS.n605 DVSS 0.31291f
C5070 VSS.t36 DVSS 4.27073f
C5071 VSS.t21 DVSS 4.57579f
C5072 VSS.t181 DVSS 1.36257f
C5073 VSS.t227 DVSS 4.16905f
C5074 VSS.t185 DVSS 4.61646f
C5075 VSS.n606 DVSS 0.671115f
C5076 VSS.t26 DVSS 0.732126f
C5077 VSS.n607 DVSS 4.57579f
C5078 VSS.n608 DVSS 0.317213f
C5079 VSS.n609 DVSS 0.201105f
C5080 VSS.n610 DVSS 0.456818f
C5081 VSS.n611 DVSS 0.154979f
C5082 VSS.n612 DVSS 0.184271f
C5083 VSS.n613 DVSS 0.184271f
C5084 VSS.t95 DVSS 4.37242f
C5085 VSS.n614 DVSS 1.64728f
C5086 VSS.t2 DVSS 2.48109f
C5087 VSS.t92 DVSS 3.43692f
C5088 VSS.n615 DVSS 0.210354f
C5089 VSS.n616 DVSS 0.210354f
C5090 VSS.n617 DVSS 0.246725f
C5091 VSS.n618 DVSS 0.053941f
C5092 VSS.n619 DVSS 0.055762f
C5093 VSS.n620 DVSS 0.324725f
C5094 VSS.t12 DVSS 4.75882f
C5095 VSS.t156 DVSS 2.11503f
C5096 VSS.n621 DVSS 0.409292f
C5097 VSS.n622 DVSS 0.404475f
C5098 VSS.n623 DVSS 0.404475f
C5099 VSS.n624 DVSS 0.898433f
C5100 VSS.t246 DVSS 5.2469f
C5101 VSS.t202 DVSS 4.75882f
C5102 VSS.t25 DVSS 5.2469f
C5103 VSS.t111 DVSS 4.75882f
C5104 VSS.t66 DVSS 5.2469f
C5105 VSS.t11 DVSS 4.75882f
C5106 VSS.t144 DVSS 5.22656f
C5107 VSS.n625 DVSS 3.82332f
C5108 VSS.n626 DVSS 0.404475f
C5109 VSS.n627 DVSS 0.404475f
C5110 VSS.n628 DVSS 0.616976f
C5111 VSS.n629 DVSS 0.898433f
C5112 VSS.n630 DVSS 0.378845f
C5113 VSS.n631 DVSS 1.22275f
C5114 VSS.n632 DVSS 0.971718f
C5115 VSS.n633 DVSS 0.971718f
C5116 VSS.n634 DVSS 0.971718f
C5117 VSS.n635 DVSS 0.971718f
C5118 VSS.n636 DVSS 0.367012f
C5119 VSS.n637 DVSS 0.129985f
C5120 VSS.n638 DVSS 1.06942f
C5121 VSS.n639 DVSS 0.1878f
C5122 VSS.n640 DVSS 0.191426f
C5123 VSS.n641 DVSS 0.862405f
C5124 VSS.n642 DVSS 0.136864f
C5125 VSS.n643 DVSS 0.135673f
C5126 VSS.n644 DVSS 0.659377f
C5127 VSS.n645 DVSS 0.649633f
C5128 VSS.n646 DVSS 0.427512f
C5129 VSS.n647 DVSS 0.427512f
C5130 VSS.n648 DVSS 0.427512f
C5131 VSS.n649 DVSS 0.427512f
C5132 VSS.n650 DVSS 0.36621f
C5133 VSS.n651 DVSS 0.089974f
C5134 VSS.n652 DVSS 0.902438f
C5135 VSS.n653 DVSS 0.594373f
C5136 VSS.n654 DVSS 0.594373f
C5137 VSS.n655 DVSS 0.594373f
C5138 VSS.n656 DVSS 0.586221f
C5139 VSS.n657 DVSS 0.035444f
C5140 VSS.n658 DVSS 0.567081f
C5141 VSS.n659 DVSS 0.594373f
C5142 VSS.n660 DVSS 0.594373f
C5143 VSS.n661 DVSS 0.594373f
C5144 VSS.n662 DVSS 0.594373f
C5145 VSS.n663 DVSS 0.680857f
C5146 VSS.n664 DVSS 0.62859f
C5147 VSS.n665 DVSS 0.20919f
C5148 VSS.n666 DVSS 0.409292f
C5149 VSS.n667 DVSS 9.80235f
C5150 VSS.n668 DVSS 0.409292f
C5151 VSS.n669 DVSS 0.698604f
C5152 VSS.n670 DVSS 1.55686f
C5153 VSS.n671 DVSS 0.136864f
C5154 VSS.n672 DVSS 0.12758f
C5155 VSS.n673 DVSS 0.139473f
C5156 VSS.n674 DVSS 0.131959f
C5157 VSS.n675 DVSS 0.176165f
C5158 VSS.n676 DVSS 0.131959f
C5159 VSS.n677 DVSS 0.03464f
C5160 VSS.n678 DVSS 0.093231f
C5161 VSS.n679 DVSS 0.145623f
C5162 VSS.n680 DVSS 0.093231f
C5163 VSS.n681 DVSS 0.187252f
C5164 VSS.n682 DVSS 0.37464f
C5165 VSS.n683 DVSS 0.285823f
C5166 VSS.n684 DVSS 0.495704f
C5167 VSS.n685 DVSS 0.450426f
C5168 VSS.n686 DVSS 0.737235f
C5169 VSS.n687 DVSS 0.779632f
C5170 VSS.n688 DVSS 1.14874f
C5171 VSS.n689 DVSS 0.122604f
C5172 VSS.n690 DVSS 0.135668f
C5173 VSS.n691 DVSS 0.409292f
C5174 VSS.n692 DVSS 2.27772f
C5175 VSS.n693 DVSS 5.34859f
C5176 VSS.n694 DVSS 0.074079f
C5177 VSS.n695 DVSS 0.376118f
C5178 VSS.n696 DVSS 0.369019f
C5179 VSS.t233 DVSS 2.78615f
C5180 VSS.t125 DVSS 4.65713f
C5181 VSS.t190 DVSS 2.78615f
C5182 VSS.n697 DVSS 0.178319f
C5183 VSS.n698 DVSS 0.178407f
C5184 VSS.n699 DVSS 0.981055f
C5185 VSS.t214 DVSS 0.506969f
C5186 VSS.n700 DVSS 1.6765f
C5187 VSS.t83 DVSS 0.412654f
C5188 VSS.n701 DVSS 1.02936f
C5189 VSS.n702 DVSS 0.294032f
C5190 VSS.n703 DVSS 5.4272f
C5191 VSS.n704 DVSS 5.71627f
C5192 VSS.t212 DVSS 0.412654f
C5193 VSS.n705 DVSS 1.02936f
C5194 VSS.t176 DVSS 0.412654f
C5195 VSS.n706 DVSS 0.253124f
C5196 VSS.n707 DVSS 0.370974f
C5197 VSS.n708 DVSS 0.201105f
C5198 VSS.n709 DVSS 0.200927f
C5199 VSS.t175 DVSS 2.23705f
C5200 VSS.t193 DVSS 2.19638f
C5201 VSS.t128 DVSS 3.29457f
C5202 VSS.t225 DVSS 1.22021f
C5203 VSS.n710 DVSS 0.094511f
C5204 VSS.n711 DVSS 0.094511f
C5205 VSS.n712 DVSS 0.616198f
C5206 VSS.n713 DVSS 0.31291f
C5207 VSS.t229 DVSS 3.92501f
C5208 VSS.t191 DVSS 2.23705f
C5209 VSS.t10 DVSS 1.56594f
C5210 VSS.n714 DVSS 3.92501f
C5211 VSS.t230 DVSS 4.51478f
C5212 VSS.t187 DVSS 1.66762f
C5213 VSS.n715 DVSS 0.080615f
C5214 VSS.n716 DVSS 0.456818f
C5215 VSS.n717 DVSS 0.398407f
C5216 VSS.n718 DVSS 0.246725f
C5217 VSS.n719 DVSS 0.391577f
C5218 VSS.n720 DVSS 0.324725f
C5219 VSS.n721 DVSS 0.210354f
C5220 VSS.t140 DVSS 0.915157f
C5221 VSS.n722 DVSS 4.00636f
C5222 VSS.n723 DVSS 0.210354f
C5223 VSS.n724 DVSS 0.053941f
C5224 VSS.n725 DVSS 0.212638f
C5225 VSS.n726 DVSS 0.737969f
C5226 VSS.n727 DVSS 0.324725f
C5227 VSS.n728 DVSS 0.210893f
C5228 VSS.n729 DVSS 3.98602f
C5229 VSS.n730 DVSS 0.335946f
C5230 VSS.n731 DVSS 2.7048f
C5231 VSS.t53 DVSS 2.35907f
C5232 VSS.t101 DVSS 4.18939f
C5233 VSS.t52 DVSS 1.56594f
C5234 VSS.n732 DVSS 0.074079f
C5235 VSS.n733 DVSS 0.376118f
C5236 VSS.n734 DVSS 0.376118f
C5237 VSS.n735 DVSS 1.70829f
C5238 VSS.n736 DVSS 0.169394f
C5239 VSS.n737 DVSS 1.6765f
C5240 VSS.n738 DVSS 0.169394f
C5241 VSS.n739 DVSS 0.169394f
C5242 VSS.n740 DVSS 0.114351f
C5243 VSS.n741 DVSS 0.153316f
C5244 VSS.n742 DVSS 0.212563f
C5245 VSS.n743 DVSS 0.212563f
C5246 VSS.n744 DVSS 0.277011f
C5247 VSS.n745 DVSS 0.277011f
C5248 VSS.n746 DVSS 0.277011f
C5249 VSS.n747 DVSS 0.277011f
C5250 VSS.n748 DVSS 0.467183f
C5251 VSS.n749 DVSS 0.139473f
C5252 VSS.n750 DVSS 0.141038f
C5253 VSS.n751 DVSS 0.523029f
C5254 VSS.n752 DVSS 0.100962f
C5255 VSS.n753 DVSS 0.256348f
C5256 VSS.n754 DVSS 0.407741f
C5257 VSS.n755 DVSS 0.211575f
C5258 VSS.n756 DVSS 0.211575f
C5259 VSS.n757 DVSS 0.211575f
C5260 VSS.n758 DVSS 0.211575f
C5261 VSS.n759 DVSS 0.184283f
C5262 VSS.n760 DVSS 0.088594f
C5263 VSS.n761 DVSS 0.011519f
C5264 VSS.n762 DVSS 0.210893f
C5265 VSS.n763 DVSS 3.80299f
C5266 VSS.n764 DVSS 1.46425f
C5267 VSS.t121 DVSS 2.23705f
C5268 VSS.n765 DVSS 1.5456f
C5269 VSS.n766 DVSS 0.096637f
C5270 VSS.t195 DVSS 2.37941f
C5271 VSS.t80 DVSS 3.0912f
C5272 VSS.n767 DVSS 4.75882f
C5273 VSS.t45 DVSS 2.1557f
C5274 VSS.t87 DVSS 0.671115f
C5275 VSS.n768 DVSS 4.41309f
C5276 VSS.t37 DVSS 4.6368f
C5277 VSS.n769 DVSS 0.094511f
C5278 VSS.t93 DVSS 0.83381f
C5279 VSS.n770 DVSS 0.094511f
C5280 VSS.n771 DVSS 0.059383f
C5281 VSS.n772 DVSS 0.406861f
C5282 VSS.n773 DVSS 0.238033f
C5283 VSS.n774 DVSS 0.067257f
C5284 VSS.n775 DVSS 0.114351f
C5285 VSS.n776 DVSS 0.059383f
C5286 VSS.n777 DVSS 0.406861f
C5287 VSS.n778 DVSS 0.238033f
C5288 VSS.n779 DVSS 0.067257f
C5289 VSS.n780 DVSS 0.114351f
C5290 VSS.n781 DVSS 0.391577f
C5291 VSS.n782 DVSS 0.616198f
C5292 VSS.n783 DVSS 0.256757f
C5293 VSS.n784 DVSS 0.132568f
C5294 VSS.n785 DVSS 0.200927f
C5295 VSS.t166 DVSS 0.412654f
C5296 VSS.n786 DVSS 1.02936f
C5297 VSS.n787 DVSS 0.294032f
C5298 VSS.t17 DVSS 0.412654f
C5299 VSS.n788 DVSS 0.31291f
C5300 VSS.t221 DVSS 2.25739f
C5301 VSS.t168 DVSS 0.506969f
C5302 VSS.n789 DVSS 3.66063f
C5303 VSS.n790 DVSS 3.96568f
C5304 VSS.t220 DVSS 0.711789f
C5305 VSS.n791 DVSS 3.06965f
C5306 VSS.n792 DVSS 0.188923f
C5307 VSS.n793 DVSS 3.57662f
C5308 VSS.n794 DVSS 2.27772f
C5309 VSS.n795 DVSS 0.369019f
C5310 VSS.n796 DVSS 1.54772f
C5311 VSS.n797 DVSS 0.949994f
C5312 VSS.n798 DVSS 0.981055f
C5313 VSS.n799 DVSS 0.080615f
C5314 VSS.n800 DVSS 0.178319f
C5315 VSS.t16 DVSS 0.142358f
C5316 VSS.n801 DVSS 0.178407f
C5317 VSS.n802 DVSS 0.253124f
C5318 VSS.n803 DVSS 0.370974f
C5319 VSS.n804 DVSS 1.2573f
C5320 VSS.n805 DVSS 0.317213f
C5321 VSS.n806 DVSS 0.752463f
C5322 VSS.n807 DVSS 2.25739f
C5323 VSS.n808 DVSS 0.096637f
C5324 VSS.n809 DVSS 0.094511f
C5325 VSS.n810 DVSS 0.153316f
C5326 VSS.n811 DVSS 1.52526f
C5327 VSS.t232 DVSS 0.305052f
C5328 VSS.n812 DVSS 3.23356f
C5329 VSS.n813 DVSS 0.096637f
C5330 VSS.n814 DVSS 0.094511f
C5331 VSS.n815 DVSS 0.059383f
C5332 VSS.n816 DVSS 0.406861f
C5333 VSS.n817 DVSS 0.238033f
C5334 VSS.n818 DVSS 0.067257f
C5335 VSS.n819 DVSS 0.169394f
C5336 VSS.n820 DVSS 0.406861f
C5337 VSS.n821 DVSS 0.059383f
C5338 VSS.n822 DVSS 0.114351f
C5339 VSS.n823 DVSS 0.153316f
C5340 VSS.n824 DVSS 0.096637f
C5341 VSS.n825 DVSS 0.955831f
C5342 VSS.t76 DVSS 0.671115f
C5343 VSS.t209 DVSS 3.864f
C5344 VSS.t15 DVSS 1.3829f
C5345 VSS.n826 DVSS 4.75882f
C5346 VSS.n827 DVSS 0.369019f
C5347 VSS.n828 DVSS 0.688262f
C5348 VSS.n829 DVSS 0.763628f
C5349 VSS.n830 DVSS 0.843255f
C5350 VSS.n831 DVSS 0.135937f
C5351 VSS.n832 DVSS 0.184271f
C5352 VSS.t240 DVSS 4.2504f
C5353 VSS.n833 DVSS 0.184271f
C5354 VSS.n834 DVSS 0.094595f
C5355 VSS.n835 DVSS 0.206313f
C5356 VSS.n836 DVSS 0.055762f
C5357 VSS.n837 DVSS 0.184271f
C5358 VSS.t203 DVSS 2.07436f
C5359 VSS.n838 DVSS 0.184271f
C5360 VSS.n839 DVSS 0.154979f
C5361 VSS.n840 DVSS 0.523872f
C5362 VSS.n841 DVSS 0.079921f
C5363 VSS.n842 DVSS 0.178319f
C5364 VSS.t211 DVSS 4.41309f
C5365 VSS.n843 DVSS 0.178319f
C5366 VSS.n844 DVSS 0.256757f
C5367 VSS.n845 DVSS 0.132568f
C5368 VSS.n846 DVSS 0.096637f
C5369 VSS.n847 DVSS 1.60661f
C5370 VSS.n848 DVSS 3.88433f
C5371 VSS.n849 DVSS 0.317213f
C5372 VSS.n850 DVSS 1.2573f
C5373 VSS.n851 DVSS 0.294032f
C5374 VSS.n852 DVSS 4.9285f
C5375 VSS.n853 DVSS 5.71627f
C5376 VSS.n854 DVSS 1.54772f
C5377 VSS.n855 DVSS 0.949994f
C5378 VSS.n856 DVSS 0.31291f
C5379 VSS.n857 DVSS 4.12838f
C5380 VSS.t117 DVSS 3.08761f
C5381 VSS.t234 DVSS 1.60633f
C5382 VSS.n858 DVSS 3.64029f
C5383 VSS.t161 DVSS 4.75882f
C5384 VSS.t231 DVSS 2.19638f
C5385 VSS.t213 DVSS 3.15221f
C5386 VSS.n859 DVSS 0.376118f
C5387 VSS.n860 DVSS 0.369019f
C5388 VSS.n861 DVSS 0.688262f
C5389 VSS.n862 DVSS 0.763628f
C5390 VSS.n863 DVSS 0.843255f
C5391 VSS.n864 DVSS 0.135937f
C5392 VSS.n865 DVSS 0.184271f
C5393 VSS.t96 DVSS 3.7013f
C5394 VSS.n866 DVSS 0.184271f
C5395 VSS.n867 DVSS 0.094595f
C5396 VSS.n868 DVSS 0.206313f
C5397 VSS.n869 DVSS 0.212638f
C5398 VSS.n870 DVSS 0.335946f
C5399 VSS.n871 DVSS 2.13537f
C5400 VSS.t186 DVSS 4.43343f
C5401 VSS.t56 DVSS 3.53861f
C5402 VSS.t239 DVSS 1.62695f
C5403 VSS.t228 DVSS 1.70829f
C5404 VSS.t97 DVSS 3.13187f
C5405 VSS.t198 DVSS 3.64029f
C5406 VSS.n872 DVSS 3.11153f
C5407 VSS.n873 DVSS 0.324725f
C5408 VSS.n874 DVSS 0.391577f
C5409 VSS.n875 DVSS 0.398407f
C5410 VSS.n876 DVSS 0.523872f
C5411 VSS.n877 DVSS 0.079921f
C5412 VSS.n878 DVSS 0.178319f
C5413 VSS.t82 DVSS 1.1592f
C5414 VSS.n879 DVSS 0.178319f
C5415 VSS.n880 DVSS 0.256757f
C5416 VSS.n881 DVSS 0.132568f
C5417 VSS.n882 DVSS 0.370974f
C5418 VSS.n883 DVSS 0.253124f
C5419 VSS.n884 DVSS 0.178407f
C5420 VSS.t22 DVSS 4.16905f
C5421 VSS.n885 DVSS 0.793136f
C5422 VSS.t33 DVSS 3.57928f
C5423 VSS.t113 DVSS 2.62345f
C5424 VSS.t1 DVSS 1.7693f
C5425 VSS.n886 DVSS 4.45377f
C5426 VSS.n887 DVSS 0.31291f
C5427 VSS.n888 DVSS 0.949994f
C5428 VSS.n889 DVSS 0.981055f
C5429 VSS.n890 DVSS 0.196483f
C5430 VSS.n891 DVSS 0.376118f
C5431 VSS.t109 DVSS 1.28122f
C5432 VSS.t20 DVSS 3.57928f
C5433 VSS.t148 DVSS 4.88084f
C5434 VSS.n892 DVSS 8.89084f
C5435 VSS.t62 DVSS 7.299661f
C5436 VSS.t63 DVSS 7.30124f
C5437 VSS.t177 DVSS 7.30124f
C5438 VSS.t137 DVSS 7.30124f
C5439 VSS.t114 DVSS 7.30124f
C5440 VSS.t38 DVSS 7.30124f
C5441 VSS.t217 DVSS 7.30124f
C5442 VSS.t24 DVSS 7.30124f
C5443 VSS.t180 DVSS 7.30124f
C5444 VSS.t107 DVSS 7.30124f
C5445 VSS.t142 DVSS 7.30124f
C5446 VSS.t94 DVSS 7.30124f
C5447 VSS.t59 DVSS 7.30124f
C5448 VSS.t7 DVSS 7.30124f
C5449 VSS.t152 DVSS 7.30124f
C5450 VSS.t131 DVSS 7.30124f
C5451 VSS.t64 DVSS 7.30124f
C5452 VSS.t61 DVSS 7.30124f
C5453 VSS.t14 DVSS 7.30124f
C5454 VSS.t98 DVSS 7.30124f
C5455 VSS.t178 DVSS 7.30124f
C5456 VSS.t85 DVSS 7.30124f
C5457 VSS.t5 DVSS 7.30124f
C5458 VSS.t35 DVSS 7.30124f
C5459 VSS.t44 DVSS 7.30124f
C5460 VSS.t65 DVSS 7.30124f
C5461 VSS.t158 DVSS 7.30124f
C5462 VSS.t170 DVSS 7.30124f
C5463 VSS.t100 DVSS 7.30124f
C5464 VSS.t164 DVSS 4.00944f
C5465 VSS.n893 DVSS 10.512199f
C5466 VSS.t132 DVSS 6.13117f
C5467 VSS.n894 DVSS 0.512107f
C5468 VSS.n895 DVSS 31.763498f
C5469 VSS.n896 DVSS 0.512107f
C5470 VSS.n897 DVSS 0.044987f
C5471 VSS.n898 DVSS 4.24715f
C5472 VSS.n899 DVSS 4.26694f
C5473 VSS.n900 DVSS 4.31057f
C5474 VSS.n901 DVSS 4.38636f
C5475 VSS.n902 DVSS 1.40198f
C5476 VSS.n903 DVSS 2.17796f
C5477 VSS.n904 DVSS 0.700166f
C5478 VSS.n905 DVSS 3.65062f
C5479 VSS.n906 DVSS 0.700166f
C5480 VSS.n907 DVSS 1.19171f
C5481 VSS.n908 DVSS 0.886472f
C5482 VSS.n909 DVSS 4.39124f
C5483 VSS.n910 DVSS 4.28957f
C5484 VSS.n911 DVSS 4.26708f
C5485 VSS.n912 DVSS 4.26654f
C5486 VSS.n913 DVSS 0.044987f
C5487 VSS.n914 DVSS 0.512107f
C5488 VSS.n915 DVSS 14.716499f
C5489 VSS.n916 DVSS 0.512107f
C5490 VSS.n917 DVSS 0.089429f
C5491 VSS.n918 DVSS 4.26317f
C5492 VSS.n919 DVSS 4.31057f
C5493 VSS.n920 DVSS 5.49314f
C5494 VSS.n921 DVSS 4.36412f
C5495 VSS.n922 DVSS 2.66264f
C5496 VSS.n923 DVSS 2.08425f
C5497 VSS.n924 DVSS 0.198295f
C5498 VSS.n925 DVSS 0.953796f
C5499 VSS.n926 DVSS 0.802851f
C5500 VSS.n927 DVSS 0.427512f
C5501 VSS.n928 DVSS 0.594373f
C5502 VSS.n929 DVSS 0.427512f
C5503 VSS.n930 DVSS 0.594373f
C5504 VSS.n931 DVSS 0.427512f
C5505 VSS.n932 DVSS 0.594373f
C5506 VSS.n933 DVSS 0.427512f
C5507 VSS.n934 DVSS 0.035444f
C5508 VSS.n935 DVSS 0.567081f
C5509 VSS.n936 DVSS 0.594373f
C5510 VSS.n937 DVSS 0.971718f
C5511 VSS.n938 DVSS 0.971718f
C5512 VSS.n939 DVSS 0.971718f
C5513 VSS.n940 DVSS 0.971718f
C5514 VSS.n941 DVSS 1.1935f
C5515 VSS.n942 DVSS 0.813153f
C5516 VSS.n943 DVSS 0.671089f
C5517 VSS.n944 DVSS 0.341792f
C5518 VSS.n945 DVSS 1.26088f
C5519 VSS.n946 DVSS 0.341792f
C5520 VSS.n947 DVSS 0.597705f
C5521 VSS.n948 DVSS 0.999855f
C5522 VSS.n949 DVSS 1.28393f
C5523 VSS.n950 DVSS 0.704567f
C5524 VSS.n951 DVSS 0.427512f
C5525 VSS.n952 DVSS 0.427512f
C5526 VSS.n953 DVSS 0.427512f
C5527 VSS.n954 DVSS 0.401638f
C5528 VSS.n955 DVSS 0.261333f
C5529 VSS.n956 DVSS 0.277011f
C5530 VSS.n957 DVSS 0.277011f
C5531 VSS.n958 DVSS 0.505013f
C5532 VSS.n959 DVSS 0.277011f
C5533 VSS.n960 DVSS 0.211575f
C5534 VSS.n961 DVSS 0.211575f
C5535 VSS.n962 DVSS 0.211575f
C5536 VSS.n963 DVSS 0.200056f
C5537 VSS.n964 DVSS 0.088594f
C5538 VSS.n965 DVSS 0.011519f
C5539 VSS.n966 DVSS 0.184283f
C5540 VSS.n967 DVSS 0.211575f
C5541 VSS.n968 DVSS 0.211575f
C5542 VSS.n969 DVSS 0.211575f
C5543 VSS.n970 DVSS 0.211575f
C5544 VSS.n971 DVSS 0.407741f
C5545 VSS.n972 DVSS 0.256348f
C5546 VSS.n973 DVSS 0.100962f
C5547 VSS.n974 DVSS 0.593348f
C5548 VSS.n975 DVSS 0.139473f
C5549 VSS.n976 DVSS 0.141038f
C5550 VSS.n977 DVSS 0.523029f
C5551 VSS.n978 DVSS 0.467183f
C5552 VSS.n979 DVSS 0.277011f
C5553 VSS.n980 DVSS 0.277011f
C5554 VSS.n981 DVSS 0.277011f
C5555 VSS.n982 DVSS 0.277011f
C5556 VSS.n983 DVSS 0.223503f
C5557 VSS.n984 DVSS 0.022701f
C5558 VSS.n985 DVSS 0.113989f
C5559 VSS.n986 DVSS 0.223152f
C5560 VSS.n987 DVSS 0.286553f
C5561 VSS.n988 DVSS 0.286553f
C5562 VSS.n989 DVSS 0.286553f
C5563 VSS.n990 DVSS 0.286553f
C5564 VSS.n991 DVSS 0.516281f
C5565 VSS.n992 DVSS 0.576971f
C5566 VSS.n993 DVSS 0.093231f
C5567 VSS.n994 DVSS 0.03464f
C5568 VSS.n995 DVSS 0.584036f
C5569 VSS.n996 DVSS 0.176165f
C5570 VSS.n997 DVSS 0.139783f
C5571 VSS.n998 DVSS 0.145623f
C5572 VSS.n999 DVSS 0.093231f
C5573 VSS.n1000 DVSS 0.031491f
C5574 VSS.n1001 DVSS 0.031682f
C5575 VSS.n1002 DVSS 0.180466f
C5576 VSS.n1003 DVSS 3.7013f
C5577 VSS.t149 DVSS 3.27423f
C5578 VSS.n1004 DVSS 0.180466f
C5579 VSS.n1005 DVSS 0.177913f
C5580 VSS.n1006 DVSS 0.053984f
C5581 VSS.n1007 DVSS 0.185526f
C5582 VSS.n1008 DVSS 0.197943f
C5583 VSS.n1009 DVSS 0.197943f
C5584 VSS.n1010 DVSS 0.197943f
C5585 VSS.n1011 DVSS 0.375281f
C5586 VSS.n1012 DVSS 0.379809f
C5587 VSS.n1013 DVSS 0.079868f
C5588 VSS.n1014 DVSS 0.124219f
C5589 VSS.n1015 DVSS 4.6368f
C5590 VSS.n1016 DVSS 1.70829f
C5591 VSS.n1017 DVSS 2.03368f
C5592 VSS.n1018 DVSS 0.124219f
C5593 VSS.n1019 DVSS 0.081219f
C5594 VSS.n1020 DVSS 0.197114f
C5595 VSS.n1021 DVSS 0.03464f
C5596 VSS.n1022 DVSS 0.036109f
C5597 VSS.n1023 DVSS 0.379809f
C5598 VSS.n1024 DVSS 0.375281f
C5599 VSS.n1025 DVSS 0.197943f
C5600 VSS.n1026 DVSS 0.197943f
C5601 VSS.n1027 DVSS 0.197943f
C5602 VSS.n1028 DVSS 0.185526f
C5603 VSS.n1029 DVSS 0.053984f
C5604 VSS.n1030 DVSS 0.156375f
C5605 VSS.n1031 DVSS 0.016184f
C5606 VSS.n1032 DVSS 0.082547f
C5607 VSS.n1033 DVSS 0.10606f
C5608 VSS.n1034 DVSS 0.10606f
C5609 VSS.n1035 DVSS 0.10606f
C5610 VSS.n1036 DVSS 0.10606f
C5611 VSS.n1037 DVSS 0.221965f
C5612 VSS.n1038 DVSS 0.112492f
C5613 VSS.n1039 DVSS 0.180466f
C5614 VSS.t106 DVSS 0.508421f
C5615 VSS.n1040 DVSS 0.180466f
C5616 VSS.n1041 DVSS 0.177913f
C5617 VSS.n1042 DVSS 0.030537f
C5618 VSS.n1043 DVSS 0.082547f
C5619 VSS.n1044 DVSS 0.10606f
C5620 VSS.n1045 DVSS 0.10606f
C5621 VSS.n1046 DVSS 0.10606f
C5622 VSS.n1047 DVSS 0.10606f
C5623 VSS.n1048 DVSS 0.180569f
C5624 VSS.n1049 DVSS 0.158957f
C5625 VSS.n1050 DVSS 0.086446f
C5626 VSS.n1051 DVSS 0.145623f
C5627 VSS.n1052 DVSS 1.99301f
C5628 VSS.n1053 DVSS 0.145623f
C5629 VSS.n1054 DVSS 0.093231f
C5630 VSS.n1055 DVSS 0.263914f
C5631 VSS.n1056 DVSS 1.42354f
C5632 VSS.n1057 DVSS 1.09633f
C5633 VSS.n1058 DVSS 0.277796f
C5634 VSS.n1059 DVSS 0.409292f
C5635 VSS.n1060 DVSS 0.122604f
C5636 VSS.n1061 DVSS 0.135668f
C5637 VSS.t86 DVSS 4.35208f
C5638 VSS.n1062 DVSS 3.15221f
C5639 VSS.t130 DVSS 2.5006f
C5640 VSS.t194 DVSS 3.1695f
C5641 VSS.t205 DVSS 0.506969f
C5642 VSS.n1063 DVSS 1.54772f
C5643 VSS.n1064 DVSS 0.369019f
C5644 VSS.n1065 DVSS 1.60661f
C5645 VSS.n1066 DVSS 4.27073f
C5646 VSS.n1067 DVSS 4.81983f
C5647 VSS.t204 DVSS 2.27772f
C5648 VSS.n1068 DVSS 0.36621f
C5649 VSS.n1069 DVSS 0.427512f
C5650 VSS.n1070 DVSS 0.545296f
C5651 VSS.n1071 DVSS 0.427512f
C5652 VSS.n1072 DVSS 0.545296f
C5653 VSS.n1073 DVSS 0.427512f
C5654 VSS.n1074 DVSS 0.545296f
C5655 VSS.n1075 DVSS 0.427512f
C5656 VSS.n1076 DVSS 0.545296f
C5657 VSS.n1077 DVSS 0.953796f
C5658 VSS.n1078 DVSS 0.697743f
C5659 VSS.n1079 DVSS 0.198295f
C5660 VSS.n1080 DVSS 0.362968f
C5661 VSS.n1081 DVSS 0.563507f
C5662 VSS.n1082 DVSS 1.1935f
C5663 VSS.n1083 DVSS 0.971718f
C5664 VSS.n1084 DVSS 0.971718f
C5665 VSS.n1085 DVSS 0.971718f
C5666 VSS.n1086 DVSS 0.971718f
C5667 VSS.n1087 DVSS 0.902438f
C5668 VSS.n1088 DVSS 0.089974f
C5669 VSS.n1089 DVSS 0.341966f
C5670 VSS.n1090 DVSS 4.90118f
C5671 VSS.n1091 DVSS 0.409292f
C5672 VSS.n1092 DVSS 0.404475f
C5673 VSS.n1093 DVSS 2.37941f
C5674 VSS.n1094 DVSS 0.404475f
C5675 VSS.n1095 DVSS 0.596772f
C5676 VSS.n1096 DVSS 0.680848f
C5677 VSS.n1097 DVSS 0.58314f
C5678 VSS.n1098 DVSS 0.545296f
C5679 VSS.n1099 DVSS 0.545296f
C5680 VSS.n1100 DVSS 0.545296f
C5681 VSS.n1101 DVSS 0.540443f
C5682 VSS.n1102 DVSS 2.54313f
C5683 VSS.n1104 DVSS 0.341966f
C5684 VSS.n1105 DVSS 3.82332f
C5685 VSS.n1106 DVSS 0.341966f
C5686 VSS.n1107 DVSS 0.341792f
C5687 VSS.n1108 DVSS 0.597705f
C5688 VSS.n1109 DVSS 0.999855f
C5689 VSS.n1110 DVSS 1.28665f
C5690 VSS.n1111 DVSS 0.974445f
C5691 VSS.n1112 DVSS 0.974445f
C5692 VSS.n1113 DVSS 0.974445f
C5693 VSS.n1114 DVSS 0.953751f
C5694 VSS.n1115 DVSS 0.089974f
C5695 VSS.n1116 DVSS 0.904756f
C5696 VSS.n1117 DVSS 0.974445f
C5697 VSS.n1118 DVSS 0.974445f
C5698 VSS.n1119 DVSS 0.974445f
C5699 VSS.n1120 DVSS 0.974445f
C5700 VSS.n1121 DVSS 1.22547f
C5701 VSS.n1122 DVSS 1.06942f
C5702 VSS.n1123 DVSS 0.191426f
C5703 VSS.n1124 DVSS 0.1878f
C5704 VSS.n1125 DVSS 0.282707f
C5705 VSS.n1126 DVSS 0.285633f
C5706 VSS.n1127 DVSS 0.135673f
C5707 VSS.n1128 DVSS 0.136864f
C5708 VSS.n1129 DVSS 0.862405f
C5709 VSS.n1130 DVSS 0.317221f
C5710 VSS.n1131 DVSS 0.255534f
C5711 VSS.n1132 DVSS 0.254689f
C5712 VSS.n1133 DVSS 4.81983f
C5713 VSS.n1134 DVSS 0.254689f
C5714 VSS.n1135 DVSS 0.255534f
C5715 VSS.n1136 DVSS 0.317221f
C5716 VSS.n1137 DVSS 0.311212f
C5717 VSS.n1138 DVSS 0.282707f
C5718 VSS.n1139 DVSS 0.285633f
C5719 VSS.n1140 DVSS 0.282707f
C5720 VSS.n1141 DVSS 0.779632f
C5721 VSS.n1142 DVSS 0.737235f
C5722 VSS.n1143 DVSS 0.450426f
C5723 VSS.n1144 DVSS 0.176165f
C5724 VSS.n1145 DVSS 2.46076f
C5725 VSS.n1146 DVSS 2.29806f
C5726 VSS.n1147 DVSS 0.145623f
C5727 VSS.n1148 DVSS 0.131959f
C5728 VSS.n1149 DVSS 0.187252f
C5729 VSS.n1150 DVSS 0.37464f
C5730 VSS.n1151 DVSS 0.285823f
C5731 VSS.n1152 DVSS 0.495704f
C5732 VSS.n1153 DVSS 0.131959f
C5733 VSS.n1154 DVSS 0.139473f
C5734 VSS.n1155 DVSS 0.593348f
C5735 VSS.n1156 DVSS 0.505013f
C5736 VSS.n1157 DVSS 0.277011f
C5737 VSS.n1158 DVSS 0.277011f
C5738 VSS.n1159 DVSS 0.277011f
C5739 VSS.n1160 DVSS 0.261333f
C5740 VSS.n1161 DVSS 0.053507f
C5741 VSS.n1162 DVSS 0.267615f
C5742 VSS.n1163 DVSS 0.286553f
C5743 VSS.n1164 DVSS 0.286553f
C5744 VSS.n1165 DVSS 0.197943f
C5745 VSS.n1166 DVSS 0.206373f
C5746 VSS.n1167 DVSS 0.197114f
C5747 VSS.n1168 DVSS 0.03464f
C5748 VSS.n1169 DVSS 0.036109f
C5749 VSS.n1170 DVSS 0.03464f
C5750 VSS.n1171 DVSS 0.031682f
C5751 VSS.n1172 DVSS 0.180466f
C5752 VSS.n1173 DVSS 0.08728f
C5753 VSS.n1174 DVSS 0.10606f
C5754 VSS.n1175 DVSS 0.10606f
C5755 VSS.n1176 DVSS 0.10606f
C5756 VSS.n1177 DVSS 0.197943f
C5757 VSS.n1178 DVSS 0.197943f
C5758 VSS.n1179 DVSS 0.185526f
C5759 VSS.n1180 DVSS 0.177913f
C5760 VSS.n1181 DVSS 0.053984f
C5761 VSS.n1182 DVSS 0.177913f
C5762 VSS.n1183 DVSS 0.180466f
C5763 VSS.n1184 DVSS 0.03485f
C5764 VSS.n1185 DVSS 0.079868f
C5765 VSS.n1186 DVSS 0.379809f
C5766 VSS.n1187 DVSS 0.375281f
C5767 VSS.n1188 DVSS 0.552922f
C5768 VSS.n1189 DVSS 0.286553f
C5769 VSS.n1190 DVSS 0.13796f
C5770 VSS.n1191 DVSS 0.13796f
C5771 VSS.n1192 DVSS 0.13796f
C5772 VSS.n1193 DVSS 0.130937f
C5773 VSS.n1194 DVSS 0.023971f
C5774 VSS.n1195 DVSS 0.022701f
C5775 VSS.n1196 DVSS 0.113989f
C5776 VSS.n1197 DVSS 0.223152f
C5777 VSS.n1198 DVSS 0.286553f
C5778 VSS.n1199 DVSS 0.286553f
C5779 VSS.n1200 DVSS 0.286553f
C5780 VSS.n1201 DVSS 0.286553f
C5781 VSS.n1202 DVSS 0.516281f
C5782 VSS.n1203 DVSS 0.576971f
C5783 VSS.n1204 DVSS 0.139783f
C5784 VSS.n1205 DVSS 0.176165f
C5785 VSS.n1206 DVSS 0.584036f
C5786 VSS.n1207 DVSS 0.03464f
C5787 VSS.n1208 DVSS 0.093231f
C5788 VSS.t146 DVSS 0.711789f
C5789 VSS.t139 DVSS 3.68097f
C5790 VSS.n1209 DVSS 4.6368f
C5791 VSS.n1210 DVSS 0.177913f
C5792 VSS.n1211 DVSS 0.08234f
C5793 VSS.n1212 DVSS 0.188923f
C5794 VSS.n1213 DVSS 5.0232f
C5795 VSS.n1214 DVSS 0.188923f
C5796 VSS.n1215 DVSS 0.191148f
C5797 VSS.n1216 DVSS 0.054985f
C5798 VSS.n1217 DVSS 0.208577f
C5799 VSS.n1218 DVSS 0.170661f
C5800 VSS.n1219 DVSS 2.37941f
C5801 VSS.n1220 DVSS 0.170661f
C5802 VSS.n1221 DVSS 0.208577f
C5803 VSS.n1222 DVSS 0.277508f
C5804 VSS.n1223 DVSS 0.13796f
C5805 VSS.n1224 DVSS 0.13796f
C5806 VSS.n1225 DVSS 0.13796f
C5807 VSS.n1226 DVSS 0.123302f
C5808 VSS.n1227 DVSS 0.075998f
C5809 VSS.n1228 DVSS 0.244293f
C5810 VSS.n1229 DVSS 0.277011f
C5811 VSS.n1230 DVSS 0.277011f
C5812 VSS.n1231 DVSS 0.505013f
C5813 VSS.n1232 DVSS 0.277011f
C5814 VSS.n1233 DVSS 0.211575f
C5815 VSS.n1234 DVSS 0.211575f
C5816 VSS.n1235 DVSS 0.211575f
C5817 VSS.n1236 DVSS 0.190663f
C5818 VSS.n1237 DVSS 0.088594f
C5819 VSS.n1238 DVSS 0.020912f
C5820 VSS.n1239 DVSS 0.184283f
C5821 VSS.n1240 DVSS 0.211575f
C5822 VSS.n1241 DVSS 0.211575f
C5823 VSS.n1242 DVSS 0.211575f
C5824 VSS.n1243 DVSS 0.211575f
C5825 VSS.n1244 DVSS 0.325199f
C5826 VSS.n1245 DVSS 0.207649f
C5827 VSS.n1246 DVSS 0.104801f
C5828 VSS.n1247 DVSS 0.240623f
C5829 VSS.n1248 DVSS 0.413161f
C5830 VSS.n1249 DVSS 0.065719f
C5831 VSS.n1250 DVSS 0.075671f
C5832 VSS.n1251 DVSS 0.096637f
C5833 VSS.n1252 DVSS 22.7431f
C5834 VSS.n1253 DVSS 0.325389f
C5835 VSS.n1254 DVSS 0.324725f
C5836 VSS.n1255 DVSS 0.184271f
C5837 VSS.n1256 DVSS 0.099748f
C5838 VSS.n1257 DVSS 0.206313f
C5839 VSS.n1258 DVSS 0.212638f
C5840 VSS.n1259 DVSS 0.335946f
C5841 VSS.n1260 DVSS 1.70829f
C5842 VSS.n1261 DVSS 1.64728f
C5843 VSS.n1262 DVSS 0.124219f
C5844 VSS.n1263 DVSS 0.081219f
C5845 VSS.n1264 DVSS 0.379809f
C5846 VSS.n1265 DVSS 0.375281f
C5847 VSS.n1266 DVSS 0.197943f
C5848 VSS.n1267 DVSS 0.10606f
C5849 VSS.n1268 DVSS 0.10606f
C5850 VSS.n1269 DVSS 0.10606f
C5851 VSS.n1270 DVSS 0.099037f
C5852 VSS.n1271 DVSS 0.030537f
C5853 VSS.n1272 DVSS 0.177913f
C5854 VSS.n1273 DVSS 5.32825f
C5855 VSS.n1274 DVSS 0.177913f
C5856 VSS.n1275 DVSS 0.01878f
C5857 VSS.n1276 DVSS 0.082547f
C5858 VSS.n1277 DVSS 0.10606f
C5859 VSS.n1278 DVSS 0.10606f
C5860 VSS.n1279 DVSS 0.10606f
C5861 VSS.n1280 DVSS 0.10606f
C5862 VSS.n1281 DVSS 0.180569f
C5863 VSS.n1282 DVSS 0.160998f
C5864 VSS.n1283 DVSS 0.10225f
C5865 VSS.n1284 DVSS 0.141147f
C5866 VSS.n1286 DVSS 0.207918f
C5867 VSS.n1287 DVSS 0.03464f
C5868 VSS.n1288 DVSS 0.093231f
C5869 VSS.t23 DVSS 0.162695f
C5870 VSS.n1289 DVSS 0.093231f
C5871 VSS.n1290 DVSS 0.163083f
C5872 VSS.n1291 DVSS 3.98058f
C5873 VSS.n1292 DVSS 6.24327f
C5874 VSS.n1293 DVSS 3.76495f
C5875 VSS.n1294 DVSS 8.33517f
C5876 VSS.n1295 DVSS 4.27708f
C5877 VSS.n1296 DVSS 0.294032f
C5878 VSS.t134 DVSS 0.412654f
C5879 VSS.n1297 DVSS 0.979944f
C5880 VSS.n1298 DVSS 0.533167f
C5881 VSS.n1299 DVSS 0.117231f
C5882 VSS.n1300 DVSS 0.178319f
C5883 VSS.t73 DVSS 2.27772f
C5884 VSS.n1301 DVSS 3.92501f
C5885 VSS.n1302 DVSS 3.53861f
C5886 VSS.n1303 DVSS 0.210893f
C5887 VSS.n1304 DVSS 0.212563f
C5888 VSS.n1305 DVSS 0.128365f
C5889 VSS.n1306 DVSS 0.341419f
C5890 VSS.n1307 DVSS 0.206767f
C5891 VSS.n1308 DVSS 2.37941f
C5892 VSS.t162 DVSS 2.62345f
C5893 VSS.t147 DVSS 2.48109f
C5894 VSS.n1309 DVSS 4.2504f
C5895 VSS.n1310 DVSS 0.369019f
C5896 VSS.n1311 DVSS 0.688262f
C5897 VSS.n1312 DVSS 0.763628f
C5898 VSS.n1313 DVSS 0.862463f
C5899 VSS.n1314 DVSS 0.135937f
C5900 VSS.n1315 DVSS 0.184271f
C5901 VSS.t90 DVSS 2.27772f
C5902 VSS.n1316 DVSS 0.184271f
C5903 VSS.n1317 DVSS 0.094595f
C5904 VSS.n1318 DVSS 0.206313f
C5905 VSS.n1319 DVSS 0.055762f
C5906 VSS.n1320 DVSS 0.184271f
C5907 VSS.t84 DVSS 3.92501f
C5908 VSS.n1321 DVSS 0.184271f
C5909 VSS.n1322 DVSS 0.154979f
C5910 VSS.n1323 DVSS 0.523872f
C5911 VSS.n1324 DVSS 0.079921f
C5912 VSS.n1325 DVSS 0.178319f
C5913 VSS.t206 DVSS 0.3864f
C5914 VSS.n1326 DVSS 0.178319f
C5915 VSS.n1327 DVSS 0.256757f
C5916 VSS.n1328 DVSS 0.132568f
C5917 VSS.n1329 DVSS 0.370974f
C5918 VSS.n1330 DVSS 0.253124f
C5919 VSS.n1331 DVSS 0.178407f
C5920 VSS.t49 DVSS 3.64029f
C5921 VSS.n1332 DVSS 0.178319f
C5922 VSS.n1333 DVSS 0.080615f
C5923 VSS.n1334 DVSS 0.981055f
C5924 VSS.n1335 DVSS 0.074079f
C5925 VSS.n1336 DVSS 0.843255f
C5926 VSS.n1337 DVSS 0.135937f
C5927 VSS.n1338 DVSS 0.184271f
C5928 VSS.t129 DVSS 2.62345f
C5929 VSS.n1339 DVSS 0.184271f
C5930 VSS.n1340 DVSS 0.094595f
C5931 VSS.n1341 DVSS 0.737969f
C5932 VSS.n1342 DVSS 0.688262f
C5933 VSS.n1343 DVSS 0.369019f
C5934 VSS.n1344 DVSS 1.64728f
C5935 VSS.t243 DVSS 4.31141f
C5936 VSS.t242 DVSS 3.3149f
C5937 VSS.n1345 DVSS 0.508421f
C5938 VSS.n1346 DVSS 0.096637f
C5939 VSS.n1347 DVSS 0.094511f
C5940 VSS.t224 DVSS 1.11853f
C5941 VSS.t19 DVSS 1.56594f
C5942 VSS.t210 DVSS 4.23006f
C5943 VSS.n1348 DVSS 4.0877f
C5944 VSS.n1349 DVSS 0.324725f
C5945 VSS.n1350 DVSS 0.391577f
C5946 VSS.n1351 DVSS 0.616198f
C5947 VSS.n1352 DVSS 0.256757f
C5948 VSS.n1353 DVSS 0.178319f
C5949 VSS.t67 DVSS 2.37941f
C5950 VSS.n1354 DVSS 0.178319f
C5951 VSS.n1355 DVSS 0.079921f
C5952 VSS.n1356 DVSS 0.456818f
C5953 VSS.t68 DVSS 0.412654f
C5954 VSS.n1357 DVSS 1.02936f
C5955 VSS.n1358 DVSS 0.294032f
C5956 VSS.n1359 DVSS 4.9285f
C5957 VSS.n1360 DVSS 5.71627f
C5958 VSS.n1361 DVSS 1.54772f
C5959 VSS.n1362 DVSS 0.369019f
C5960 VSS.n1363 DVSS 2.98951f
C5961 VSS.t46 DVSS 4.8605f
C5962 VSS.t244 DVSS 2.74547f
C5963 VSS.t69 DVSS 2.50143f
C5964 VSS.t236 DVSS 4.75882f
C5965 VSS.t222 DVSS 3.33524f
C5966 VSS.n1364 DVSS 2.01335f
C5967 VSS.n1365 DVSS 0.369019f
C5968 VSS.n1366 DVSS 0.688262f
C5969 VSS.n1367 DVSS 0.763628f
C5970 VSS.n1368 DVSS 0.843255f
C5971 VSS.n1369 DVSS 0.135937f
C5972 VSS.n1370 DVSS 0.184271f
C5973 VSS.t201 DVSS 5.71465f
C5974 VSS.n1371 DVSS 0.184271f
C5975 VSS.n1372 DVSS 0.094595f
C5976 VSS.n1373 DVSS 0.206313f
C5977 VSS.n1374 DVSS 0.055762f
C5978 VSS.n1375 DVSS 0.184271f
C5979 VSS.t78 DVSS 3.55895f
C5980 VSS.n1376 DVSS 0.184271f
C5981 VSS.n1377 DVSS 0.154979f
C5982 VSS.n1378 DVSS 0.523872f
C5983 VSS.n1379 DVSS 0.079921f
C5984 VSS.n1380 DVSS 0.178319f
C5985 VSS.t165 DVSS 3.68097f
C5986 VSS.n1381 DVSS 3.27423f
C5987 VSS.n1382 DVSS 0.177913f
C5988 VSS.n1383 DVSS 0.08234f
C5989 VSS.n1384 DVSS 0.188923f
C5990 VSS.n1385 DVSS 5.20623f
C5991 VSS.n1386 DVSS 0.188923f
C5992 VSS.n1387 DVSS 0.191148f
C5993 VSS.n1388 DVSS 0.054985f
C5994 VSS.n1389 DVSS 0.208577f
C5995 VSS.n1390 DVSS 0.170661f
C5996 VSS.n1391 DVSS 2.37941f
C5997 VSS.n1392 DVSS 0.170661f
C5998 VSS.n1393 DVSS 0.208577f
C5999 VSS.n1394 DVSS 0.277508f
C6000 VSS.n1395 DVSS 0.13796f
C6001 VSS.n1396 DVSS 0.13796f
C6002 VSS.n1397 DVSS 0.13796f
C6003 VSS.n1398 DVSS 0.123302f
C6004 VSS.n1399 DVSS 0.075998f
C6005 VSS.n1400 DVSS 0.713128f
C6006 VSS.n1401 DVSS 0.210893f
C6007 VSS.n1402 DVSS 3.96568f
C6008 VSS.n1403 DVSS 0.210893f
C6009 VSS.n1404 DVSS 0.212563f
C6010 VSS.n1405 DVSS 0.128365f
C6011 VSS.n1406 DVSS 0.341419f
C6012 VSS.n1407 DVSS 0.206767f
C6013 VSS.n1408 DVSS 2.37941f
C6014 VSS.n1409 DVSS 0.206767f
C6015 VSS.n1410 DVSS 0.341419f
C6016 VSS.n1411 DVSS 0.421535f
C6017 VSS.n1412 DVSS 0.211575f
C6018 VSS.n1413 DVSS 0.211575f
C6019 VSS.n1414 DVSS 0.211575f
C6020 VSS.n1415 DVSS 0.190663f
C6021 VSS.n1416 DVSS 0.088594f
C6022 VSS.n1417 DVSS 0.046972f
C6023 VSS.n1418 DVSS 0.254689f
C6024 VSS.n1419 DVSS 4.43343f
C6025 VSS.n1420 DVSS 0.254689f
C6026 VSS.n1421 DVSS 0.255534f
C6027 VSS.n1422 DVSS 0.317221f
C6028 VSS.n1423 DVSS 0.311212f
C6029 VSS.n1424 DVSS 0.282707f
C6030 VSS.n1425 DVSS 2.37941f
C6031 VSS.n1426 DVSS 0.282707f
C6032 VSS.n1427 DVSS 0.311212f
C6033 VSS.n1428 DVSS 0.518818f
C6034 VSS.n1429 DVSS 0.999855f
C6035 VSS.n1430 DVSS 1.28393f
C6036 VSS.n1431 DVSS 0.971718f
C6037 VSS.n1432 DVSS 0.971718f
C6038 VSS.n1433 DVSS 0.971718f
C6039 VSS.n1434 DVSS 0.951024f
C6040 VSS.n1435 DVSS 0.089974f
C6041 VSS.n1436 DVSS 0.254689f
C6042 VSS.n1437 DVSS 4.51478f
C6043 VSS.n1438 DVSS 3.74198f
C6044 VSS.n1439 DVSS 0.096637f
C6045 VSS.n1440 DVSS 0.153316f
C6046 VSS.n1441 DVSS 0.235252f
C6047 VSS.n1442 DVSS 0.066582f
C6048 x9.V2.t70 DVSS 1.00605f
C6049 x9.V2.t54 DVSS 0.105694f
C6050 x9.V2.t55 DVSS 0.105694f
C6051 x9.V2.n0 DVSS 0.215568f
C6052 x9.V2.n1 DVSS 0.425847f
C6053 x9.V2.n2 DVSS 0.133159f
C6054 x9.V2.n3 DVSS 0.192547f
C6055 x9.V2.t57 DVSS 0.031737f
C6056 x9.V2.n4 DVSS 0.152499f
C6057 x9.V2.t7 DVSS 0.031737f
C6058 x9.V2.n5 DVSS 0.140724f
C6059 x9.V2.t24 DVSS 0.031737f
C6060 x9.V2.n6 DVSS 0.140724f
C6061 x9.V2.t4 DVSS 0.031737f
C6062 x9.V2.n7 DVSS 0.140724f
C6063 x9.V2.t31 DVSS 0.031737f
C6064 x9.V2.n8 DVSS 0.140724f
C6065 x9.V2.t25 DVSS 0.031737f
C6066 x9.V2.n9 DVSS 0.140724f
C6067 x9.V2.t46 DVSS 0.031737f
C6068 x9.V2.n10 DVSS 0.140724f
C6069 x9.V2.t2 DVSS 0.031737f
C6070 x9.V2.n11 DVSS 0.140724f
C6071 x9.V2.t15 DVSS 0.031737f
C6072 x9.V2.n12 DVSS 0.140724f
C6073 x9.V2.t65 DVSS 0.031737f
C6074 x9.V2.n13 DVSS 0.140724f
C6075 x9.V2.t53 DVSS 0.031737f
C6076 x9.V2.n14 DVSS 0.140724f
C6077 x9.V2.t48 DVSS 0.031737f
C6078 x9.V2.n15 DVSS 0.140724f
C6079 x9.V2.t11 DVSS 0.031737f
C6080 x9.V2.n16 DVSS 0.140724f
C6081 x9.V2.t18 DVSS 0.031737f
C6082 x9.V2.n17 DVSS 0.140724f
C6083 x9.V2.t33 DVSS 0.031737f
C6084 x9.V2.n18 DVSS 0.140724f
C6085 x9.V2.t64 DVSS 0.031737f
C6086 x9.V2.n19 DVSS 0.140724f
C6087 x9.V2.t58 DVSS 0.031737f
C6088 x9.V2.n20 DVSS 0.140724f
C6089 x9.V2.t27 DVSS 0.031737f
C6090 x9.V2.n21 DVSS 0.140724f
C6091 x9.V2.t30 DVSS 0.031737f
C6092 x9.V2.n22 DVSS 0.140724f
C6093 x9.V2.t22 DVSS 0.031737f
C6094 x9.V2.n23 DVSS 0.140724f
C6095 x9.V2.t14 DVSS 0.031737f
C6096 x9.V2.n24 DVSS 0.140724f
C6097 x9.V2.t39 DVSS 0.031737f
C6098 x9.V2.n25 DVSS 0.140724f
C6099 x9.V2.t40 DVSS 0.031737f
C6100 x9.V2.n26 DVSS 0.140724f
C6101 x9.V2.t37 DVSS 0.031737f
C6102 x9.V2.n27 DVSS 0.140724f
C6103 x9.V2.t42 DVSS 0.031737f
C6104 x9.V2.n28 DVSS 0.140724f
C6105 x9.V2.t21 DVSS 0.031737f
C6106 x9.V2.n29 DVSS 0.140724f
C6107 x9.V2.t20 DVSS 0.031737f
C6108 x9.V2.n30 DVSS 0.140724f
C6109 x9.V2.t0 DVSS 0.114356f
C6110 x9.V2.n31 DVSS 0.058105f
C6111 x9.V2.t36 DVSS 0.031737f
C6112 x9.V2.n32 DVSS 0.140724f
C6113 x9.V2.t26 DVSS 0.031737f
C6114 x9.V2.n33 DVSS 0.140724f
C6115 x9.V2.t66 DVSS 0.031737f
C6116 x9.V2.n34 DVSS 0.140724f
C6117 x9.V2.t1 DVSS 0.031737f
C6118 x9.V2.n35 DVSS 0.140724f
C6119 x9.V2.t69 DVSS 0.031737f
C6120 x9.V2.n36 DVSS 0.140724f
C6121 x9.V2.t29 DVSS 0.031737f
C6122 x9.V2.n37 DVSS 0.140724f
C6123 x9.V2.t8 DVSS 0.031737f
C6124 x9.V2.n38 DVSS 0.140724f
C6125 x9.V2.t35 DVSS 0.031737f
C6126 x9.V2.n39 DVSS 0.140724f
C6127 x9.V2.t51 DVSS 0.031737f
C6128 x9.V2.n40 DVSS 0.140724f
C6129 x9.V2.t23 DVSS 0.031737f
C6130 x9.V2.n41 DVSS 0.140724f
C6131 x9.V2.t68 DVSS 0.031737f
C6132 x9.V2.n42 DVSS 0.140724f
C6133 x9.V2.t47 DVSS 0.031737f
C6134 x9.V2.n43 DVSS 0.140724f
C6135 x9.V2.t63 DVSS 0.031737f
C6136 x9.V2.n44 DVSS 0.140724f
C6137 x9.V2.t67 DVSS 0.031737f
C6138 x9.V2.n45 DVSS 0.140724f
C6139 x9.V2.t56 DVSS 0.031737f
C6140 x9.V2.n46 DVSS 0.140724f
C6141 x9.V2.t19 DVSS 0.031737f
C6142 x9.V2.n47 DVSS 0.140724f
C6143 x9.V2.t10 DVSS 0.031737f
C6144 x9.V2.n48 DVSS 0.140724f
C6145 x9.V2.t34 DVSS 0.031737f
C6146 x9.V2.n49 DVSS 0.140724f
C6147 x9.V2.t6 DVSS 0.031737f
C6148 x9.V2.n50 DVSS 0.140724f
C6149 x9.V2.t41 DVSS 0.031737f
C6150 x9.V2.n51 DVSS 0.140724f
C6151 x9.V2.t16 DVSS 0.031737f
C6152 x9.V2.n52 DVSS 0.140724f
C6153 x9.V2.t62 DVSS 0.031737f
C6154 x9.V2.n53 DVSS 0.140724f
C6155 x9.V2.t43 DVSS 0.031737f
C6156 x9.V2.n54 DVSS 0.327637f
C6157 x9.V2.n55 DVSS 0.192547f
C6158 x9.V2.n56 DVSS 0.192547f
C6159 x9.V2.n57 DVSS 0.192547f
C6160 x9.V2.n58 DVSS 0.192547f
C6161 x9.V2.n59 DVSS 0.192547f
C6162 x9.V2.n60 DVSS 0.192547f
C6163 x9.V2.n61 DVSS 0.192547f
C6164 x9.V2.n62 DVSS 0.192547f
C6165 x9.V2.n63 DVSS 0.192547f
C6166 x9.V2.n64 DVSS 0.192547f
C6167 x9.V2.n65 DVSS 0.192547f
C6168 x9.V2.n66 DVSS 0.192547f
C6169 x9.V2.n67 DVSS 0.192547f
C6170 x9.V2.n68 DVSS 0.192547f
C6171 x9.V2.n69 DVSS 0.192547f
C6172 x9.V2.n70 DVSS 0.192547f
C6173 x9.V2.n71 DVSS 0.192547f
C6174 x9.V2.n72 DVSS 0.192547f
C6175 x9.V2.n73 DVSS 0.192547f
C6176 x9.V2.n74 DVSS 0.192547f
C6177 x9.V2.n75 DVSS 0.192547f
C6178 x9.V2.n76 DVSS 0.192547f
C6179 x9.V2.n77 DVSS 0.192547f
C6180 x9.V2.n78 DVSS 0.192547f
C6181 x9.V2.n79 DVSS 0.192547f
C6182 x9.V2.n80 DVSS 0.192547f
C6183 x9.V2.n81 DVSS 0.192547f
C6184 x9.V2.n82 DVSS 0.192547f
C6185 x9.V2.n83 DVSS 0.192547f
C6186 x9.V2.n84 DVSS 0.192547f
C6187 x9.V2.n85 DVSS 0.192547f
C6188 x9.V2.n86 DVSS 0.192547f
C6189 x9.V2.n87 DVSS 0.192547f
C6190 x9.V2.n88 DVSS 0.192547f
C6191 x9.V2.n89 DVSS 0.192547f
C6192 x9.V2.n90 DVSS 0.192547f
C6193 x9.V2.n91 DVSS 0.192547f
C6194 x9.V2.n92 DVSS 0.192547f
C6195 x9.V2.n93 DVSS 0.192547f
C6196 x9.V2.n94 DVSS 0.192547f
C6197 x9.V2.n95 DVSS 0.192547f
C6198 x9.V2.n96 DVSS 0.192547f
C6199 x9.V2.n97 DVSS 0.192547f
C6200 x9.V2.n98 DVSS 0.192547f
C6201 x9.V2.n99 DVSS 0.192547f
C6202 x9.V2.n100 DVSS 0.192547f
C6203 x9.V2.n101 DVSS 0.192547f
C6204 x9.V2.n102 DVSS 0.192547f
C6205 x9.V2.n103 DVSS 0.192547f
C6206 x9.V2.n104 DVSS 0.140724f
C6207 x9.V2.t61 DVSS 0.031737f
C6208 x9.V2.n105 DVSS 0.140724f
C6209 x9.V2.t52 DVSS 0.031737f
C6210 x9.V2.n106 DVSS 0.140724f
C6211 x9.V2.t9 DVSS 0.031737f
C6212 x9.V2.n107 DVSS 0.140724f
C6213 x9.V2.t38 DVSS 0.031737f
C6214 x9.V2.n108 DVSS 0.140724f
C6215 x9.V2.t3 DVSS 0.031737f
C6216 x9.V2.n109 DVSS 0.140724f
C6217 x9.V2.t5 DVSS 0.031737f
C6218 x9.V2.n110 DVSS 0.140724f
C6219 x9.V2.t60 DVSS 0.031737f
C6220 x9.V2.n111 DVSS 0.140724f
C6221 x9.V2.t28 DVSS 0.031737f
C6222 x9.V2.n112 DVSS 0.140724f
C6223 x9.V2.t44 DVSS 0.031737f
C6224 x9.V2.n113 DVSS 0.140724f
C6225 x9.V2.t13 DVSS 0.031737f
C6226 x9.V2.n114 DVSS 0.140724f
C6227 x9.V2.t32 DVSS 0.031737f
C6228 x9.V2.n115 DVSS 0.140724f
C6229 x9.V2.t59 DVSS 0.031737f
C6230 x9.V2.n116 DVSS 0.192547f
C6231 x9.V2.n117 DVSS 0.192547f
C6232 x9.V2.n118 DVSS 0.192547f
C6233 x9.V2.n119 DVSS 0.192547f
C6234 x9.V2.n120 DVSS 0.192547f
C6235 x9.V2.n121 DVSS 0.192547f
C6236 x9.V2.n122 DVSS 0.192547f
C6237 x9.V2.n123 DVSS 0.192547f
C6238 x9.V2.n124 DVSS 0.329928f
C6239 x9.V2.n125 DVSS 0.152699f
C6240 x9.V2.n126 DVSS 8.880599f
C6241 x9.V2.t12 DVSS 0.031737f
C6242 x9.V2.n127 DVSS 0.140724f
C6243 x9.V2.n128 DVSS 0.154754f
C6244 x9.V2.n129 DVSS 2.44267f
C6245 x9.V2.n130 DVSS 2.90206f
C6246 x9.V2.t50 DVSS 0.105694f
C6247 x9.V2.t49 DVSS 0.105694f
C6248 x9.V2.n131 DVSS 0.215568f
C6249 x9.V2.n132 DVSS 0.411861f
C6250 x9.V2.n133 DVSS 0.437043f
C6251 x9.V2.n134 DVSS 0.156394f
C6252 x9.V2.t17 DVSS 0.223553f
C6253 x9.V2.t45 DVSS 0.369599f
C6254 x9.V2.n135 DVSS 0.837759f
C6255 x9.V2.n136 DVSS 0.859643f
C6256 x9.V2.n137 DVSS 0.467495f
C6257 x6.V1.t53 DVSS 0.135038f
C6258 x6.V1.t94 DVSS 1.41004f
C6259 x6.V1.n0 DVSS 1.00384f
C6260 x6.V1.t81 DVSS 0.044303f
C6261 x6.V1.n1 DVSS 0.199346f
C6262 x6.V1.n2 DVSS 0.26969f
C6263 x6.V1.t79 DVSS 0.044303f
C6264 x6.V1.n3 DVSS 0.214352f
C6265 x6.V1.t13 DVSS 0.044303f
C6266 x6.V1.n4 DVSS 0.196967f
C6267 x6.V1.t37 DVSS 0.044303f
C6268 x6.V1.n5 DVSS 0.196967f
C6269 x6.V1.t10 DVSS 0.044303f
C6270 x6.V1.n6 DVSS 0.196967f
C6271 x6.V1.t44 DVSS 0.044303f
C6272 x6.V1.n7 DVSS 0.196967f
C6273 x6.V1.t38 DVSS 0.044303f
C6274 x6.V1.n8 DVSS 0.196967f
C6275 x6.V1.t64 DVSS 0.044303f
C6276 x6.V1.n9 DVSS 0.196967f
C6277 x6.V1.t8 DVSS 0.044303f
C6278 x6.V1.n10 DVSS 0.196967f
C6279 x6.V1.t28 DVSS 0.044303f
C6280 x6.V1.n11 DVSS 0.196967f
C6281 x6.V1.t89 DVSS 0.044303f
C6282 x6.V1.n12 DVSS 0.196967f
C6283 x6.V1.t72 DVSS 0.044303f
C6284 x6.V1.n13 DVSS 0.196967f
C6285 x6.V1.t66 DVSS 0.044303f
C6286 x6.V1.n14 DVSS 0.196967f
C6287 x6.V1.t21 DVSS 0.044303f
C6288 x6.V1.n15 DVSS 0.196967f
C6289 x6.V1.t31 DVSS 0.044303f
C6290 x6.V1.n16 DVSS 0.196967f
C6291 x6.V1.t46 DVSS 0.044303f
C6292 x6.V1.n17 DVSS 0.196967f
C6293 x6.V1.t88 DVSS 0.044303f
C6294 x6.V1.n18 DVSS 0.196967f
C6295 x6.V1.t80 DVSS 0.044303f
C6296 x6.V1.n19 DVSS 0.196967f
C6297 x6.V1.t40 DVSS 0.044303f
C6298 x6.V1.n20 DVSS 0.196967f
C6299 x6.V1.t43 DVSS 0.044303f
C6300 x6.V1.n21 DVSS 0.196967f
C6301 x6.V1.t35 DVSS 0.044303f
C6302 x6.V1.n22 DVSS 0.196967f
C6303 x6.V1.t26 DVSS 0.044303f
C6304 x6.V1.n23 DVSS 0.196967f
C6305 x6.V1.t52 DVSS 0.044303f
C6306 x6.V1.n24 DVSS 0.196967f
C6307 x6.V1.t54 DVSS 0.044303f
C6308 x6.V1.n25 DVSS 0.196967f
C6309 x6.V1.t50 DVSS 0.044303f
C6310 x6.V1.n26 DVSS 0.196967f
C6311 x6.V1.t57 DVSS 0.044303f
C6312 x6.V1.n27 DVSS 0.196967f
C6313 x6.V1.t34 DVSS 0.044303f
C6314 x6.V1.n28 DVSS 0.196967f
C6315 x6.V1.t33 DVSS 0.044303f
C6316 x6.V1.n29 DVSS 0.196967f
C6317 x6.V1.t1 DVSS 0.044303f
C6318 x6.V1.n30 DVSS 0.196967f
C6319 x6.V1.t49 DVSS 0.044303f
C6320 x6.V1.n31 DVSS 0.196967f
C6321 x6.V1.t39 DVSS 0.044303f
C6322 x6.V1.n32 DVSS 0.196967f
C6323 x6.V1.t90 DVSS 0.044303f
C6324 x6.V1.n33 DVSS 0.196967f
C6325 x6.V1.t7 DVSS 0.044303f
C6326 x6.V1.n34 DVSS 0.196967f
C6327 x6.V1.t93 DVSS 0.044303f
C6328 x6.V1.n35 DVSS 0.196967f
C6329 x6.V1.t42 DVSS 0.044303f
C6330 x6.V1.n36 DVSS 0.196967f
C6331 x6.V1.t16 DVSS 0.044303f
C6332 x6.V1.n37 DVSS 0.196967f
C6333 x6.V1.t48 DVSS 0.044303f
C6334 x6.V1.n38 DVSS 0.196967f
C6335 x6.V1.t67 DVSS 0.044303f
C6336 x6.V1.n39 DVSS 0.196967f
C6337 x6.V1.t36 DVSS 0.044303f
C6338 x6.V1.n40 DVSS 0.196967f
C6339 x6.V1.t92 DVSS 0.044303f
C6340 x6.V1.n41 DVSS 0.196967f
C6341 x6.V1.t65 DVSS 0.044303f
C6342 x6.V1.n42 DVSS 0.196967f
C6343 x6.V1.t87 DVSS 0.044303f
C6344 x6.V1.n43 DVSS 0.196967f
C6345 x6.V1.t91 DVSS 0.044303f
C6346 x6.V1.n44 DVSS 0.196967f
C6347 x6.V1.t78 DVSS 0.044303f
C6348 x6.V1.n45 DVSS 0.196967f
C6349 x6.V1.t32 DVSS 0.044303f
C6350 x6.V1.n46 DVSS 0.196967f
C6351 x6.V1.t20 DVSS 0.044303f
C6352 x6.V1.n47 DVSS 0.196967f
C6353 x6.V1.t47 DVSS 0.044303f
C6354 x6.V1.n48 DVSS 0.196967f
C6355 x6.V1.t12 DVSS 0.044303f
C6356 x6.V1.n49 DVSS 0.196967f
C6357 x6.V1.t56 DVSS 0.044303f
C6358 x6.V1.n50 DVSS 0.196967f
C6359 x6.V1.t30 DVSS 0.044303f
C6360 x6.V1.n51 DVSS 0.196967f
C6361 x6.V1.t86 DVSS 0.044303f
C6362 x6.V1.n52 DVSS 0.196967f
C6363 x6.V1.t62 DVSS 0.044303f
C6364 x6.V1.n53 DVSS 0.196967f
C6365 x6.V1.t85 DVSS 0.044303f
C6366 x6.V1.n54 DVSS 0.196967f
C6367 x6.V1.t24 DVSS 0.044303f
C6368 x6.V1.n55 DVSS 0.196967f
C6369 x6.V1.t68 DVSS 0.044303f
C6370 x6.V1.n56 DVSS 0.196967f
C6371 x6.V1.t19 DVSS 0.044303f
C6372 x6.V1.n57 DVSS 0.196967f
C6373 x6.V1.t51 DVSS 0.044303f
C6374 x6.V1.n58 DVSS 0.196967f
C6375 x6.V1.t9 DVSS 0.044303f
C6376 x6.V1.n59 DVSS 0.196967f
C6377 x6.V1.t11 DVSS 0.044303f
C6378 x6.V1.n60 DVSS 0.196967f
C6379 x6.V1.t84 DVSS 0.044303f
C6380 x6.V1.n61 DVSS 0.196967f
C6381 x6.V1.t41 DVSS 0.044303f
C6382 x6.V1.n62 DVSS 0.196967f
C6383 x6.V1.t63 DVSS 0.044303f
C6384 x6.V1.n63 DVSS 0.469622f
C6385 x6.V1.n64 DVSS 0.26969f
C6386 x6.V1.n65 DVSS 0.26969f
C6387 x6.V1.n66 DVSS 0.26969f
C6388 x6.V1.n67 DVSS 0.26969f
C6389 x6.V1.n68 DVSS 0.26969f
C6390 x6.V1.n69 DVSS 0.26969f
C6391 x6.V1.n70 DVSS 0.26969f
C6392 x6.V1.n71 DVSS 0.26969f
C6393 x6.V1.n72 DVSS 0.26969f
C6394 x6.V1.n73 DVSS 0.26969f
C6395 x6.V1.n74 DVSS 0.26969f
C6396 x6.V1.n75 DVSS 0.26969f
C6397 x6.V1.n76 DVSS 0.26969f
C6398 x6.V1.n77 DVSS 0.26969f
C6399 x6.V1.n78 DVSS 0.26969f
C6400 x6.V1.n79 DVSS 0.26969f
C6401 x6.V1.n80 DVSS 0.26969f
C6402 x6.V1.n81 DVSS 0.26969f
C6403 x6.V1.n82 DVSS 0.26969f
C6404 x6.V1.n83 DVSS 0.26969f
C6405 x6.V1.n84 DVSS 0.26969f
C6406 x6.V1.n85 DVSS 0.26969f
C6407 x6.V1.n86 DVSS 0.26969f
C6408 x6.V1.n87 DVSS 0.26969f
C6409 x6.V1.n88 DVSS 0.26969f
C6410 x6.V1.n89 DVSS 0.26969f
C6411 x6.V1.n90 DVSS 0.26969f
C6412 x6.V1.n91 DVSS 0.26969f
C6413 x6.V1.n92 DVSS 0.26969f
C6414 x6.V1.n93 DVSS 0.26969f
C6415 x6.V1.n94 DVSS 0.26969f
C6416 x6.V1.n95 DVSS 0.26969f
C6417 x6.V1.n96 DVSS 0.26969f
C6418 x6.V1.n97 DVSS 0.26969f
C6419 x6.V1.n98 DVSS 0.26969f
C6420 x6.V1.n99 DVSS 0.26969f
C6421 x6.V1.n100 DVSS 0.26969f
C6422 x6.V1.n101 DVSS 0.26969f
C6423 x6.V1.n102 DVSS 0.26969f
C6424 x6.V1.n103 DVSS 0.26969f
C6425 x6.V1.n104 DVSS 0.26969f
C6426 x6.V1.n105 DVSS 0.26969f
C6427 x6.V1.n106 DVSS 0.26969f
C6428 x6.V1.n107 DVSS 0.26969f
C6429 x6.V1.n108 DVSS 0.26969f
C6430 x6.V1.n109 DVSS 0.26969f
C6431 x6.V1.n110 DVSS 0.26969f
C6432 x6.V1.n111 DVSS 0.26969f
C6433 x6.V1.n112 DVSS 0.26969f
C6434 x6.V1.n113 DVSS 0.26969f
C6435 x6.V1.n114 DVSS 0.26969f
C6436 x6.V1.n115 DVSS 0.26969f
C6437 x6.V1.n116 DVSS 0.26969f
C6438 x6.V1.n117 DVSS 0.26969f
C6439 x6.V1.n118 DVSS 0.26969f
C6440 x6.V1.n119 DVSS 0.26969f
C6441 x6.V1.n120 DVSS 0.26969f
C6442 x6.V1.n121 DVSS 0.26969f
C6443 x6.V1.n122 DVSS 0.26969f
C6444 x6.V1.n123 DVSS 0.196967f
C6445 x6.V1.t25 DVSS 0.044303f
C6446 x6.V1.n124 DVSS 0.196967f
C6447 x6.V1.n125 DVSS 12.455999f
C6448 x6.V1.t45 DVSS 0.044303f
C6449 x6.V1.n126 DVSS 0.196967f
C6450 x6.V1.n127 DVSS 0.234774f
C6451 x6.V1.n128 DVSS 2.50125f
C6452 x6.V1.n129 DVSS 10.2707f
C6453 x6.V1.t2 DVSS 0.034299f
C6454 x6.V1.t27 DVSS 0.034299f
C6455 x6.V1.n130 DVSS 0.106673f
C6456 x6.V1.n131 DVSS 2.60019f
C6457 x6.V1.t61 DVSS 0.034299f
C6458 x6.V1.t18 DVSS 0.034299f
C6459 x6.V1.n132 DVSS 0.106673f
C6460 x6.V1.n133 DVSS 0.201325f
C6461 x6.V1.t23 DVSS 0.034299f
C6462 x6.V1.t5 DVSS 0.034299f
C6463 x6.V1.n134 DVSS 0.106673f
C6464 x6.V1.n135 DVSS 0.201325f
C6465 x6.V1.t6 DVSS 0.034299f
C6466 x6.V1.t70 DVSS 0.034299f
C6467 x6.V1.n136 DVSS 0.106673f
C6468 x6.V1.n137 DVSS 0.201325f
C6469 x6.V1.t71 DVSS 0.034299f
C6470 x6.V1.t4 DVSS 0.034299f
C6471 x6.V1.n138 DVSS 0.106673f
C6472 x6.V1.n139 DVSS 0.201228f
C6473 x6.V1.t0 DVSS 0.034299f
C6474 x6.V1.t22 DVSS 0.034299f
C6475 x6.V1.n140 DVSS 0.106673f
C6476 x6.V1.n141 DVSS 0.201228f
C6477 x6.V1.t55 DVSS 0.034299f
C6478 x6.V1.t3 DVSS 0.034299f
C6479 x6.V1.n142 DVSS 0.106673f
C6480 x6.V1.n143 DVSS 0.238096f
C6481 x6.V1.t76 DVSS 0.034143f
C6482 x6.V1.t74 DVSS 0.034143f
C6483 x6.V1.n144 DVSS 0.106107f
C6484 x6.V1.n145 DVSS 0.237588f
C6485 x6.V1.t77 DVSS 0.034143f
C6486 x6.V1.t58 DVSS 0.034143f
C6487 x6.V1.n146 DVSS 0.106107f
C6488 x6.V1.n147 DVSS 0.20072f
C6489 x6.V1.t60 DVSS 0.034143f
C6490 x6.V1.t75 DVSS 0.034143f
C6491 x6.V1.n148 DVSS 0.106107f
C6492 x6.V1.n149 DVSS 0.20072f
C6493 x6.V1.t73 DVSS 0.034143f
C6494 x6.V1.t59 DVSS 0.034143f
C6495 x6.V1.n150 DVSS 0.106107f
C6496 x6.V1.n151 DVSS 0.237588f
C6497 x6.V1.t15 DVSS 0.036247f
C6498 x6.V1.t14 DVSS 0.036247f
C6499 x6.V1.n152 DVSS 0.113646f
C6500 x6.V1.n153 DVSS 0.245774f
C6501 x6.V1.t17 DVSS 0.036247f
C6502 x6.V1.t83 DVSS 0.036247f
C6503 x6.V1.n154 DVSS 0.113646f
C6504 x6.V1.n155 DVSS 0.245774f
C6505 x6.V1.t82 DVSS 0.037962f
C6506 x6.V1.t69 DVSS 0.037962f
C6507 x6.V1.n156 DVSS 0.122278f
C6508 x6.V1.n157 DVSS 0.286804f
C6509 x6.V1.t29 DVSS 0.16958f
C6510 x6.V1.n158 DVSS 0.319705f
C6511 x6.V1.n159 DVSS 0.210087f
.ends

