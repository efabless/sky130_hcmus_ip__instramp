magic
tech sky130A
magscale 1 2
timestamp 1717127688
<< pwell >>
rect -2005 -698 2005 698
<< mvnmos >>
rect -1777 -440 -1577 440
rect -1519 -440 -1319 440
rect -1261 -440 -1061 440
rect -1003 -440 -803 440
rect -745 -440 -545 440
rect -487 -440 -287 440
rect -229 -440 -29 440
rect 29 -440 229 440
rect 287 -440 487 440
rect 545 -440 745 440
rect 803 -440 1003 440
rect 1061 -440 1261 440
rect 1319 -440 1519 440
rect 1577 -440 1777 440
<< mvndiff >>
rect -1835 428 -1777 440
rect -1835 -428 -1823 428
rect -1789 -428 -1777 428
rect -1835 -440 -1777 -428
rect -1577 428 -1519 440
rect -1577 -428 -1565 428
rect -1531 -428 -1519 428
rect -1577 -440 -1519 -428
rect -1319 428 -1261 440
rect -1319 -428 -1307 428
rect -1273 -428 -1261 428
rect -1319 -440 -1261 -428
rect -1061 428 -1003 440
rect -1061 -428 -1049 428
rect -1015 -428 -1003 428
rect -1061 -440 -1003 -428
rect -803 428 -745 440
rect -803 -428 -791 428
rect -757 -428 -745 428
rect -803 -440 -745 -428
rect -545 428 -487 440
rect -545 -428 -533 428
rect -499 -428 -487 428
rect -545 -440 -487 -428
rect -287 428 -229 440
rect -287 -428 -275 428
rect -241 -428 -229 428
rect -287 -440 -229 -428
rect -29 428 29 440
rect -29 -428 -17 428
rect 17 -428 29 428
rect -29 -440 29 -428
rect 229 428 287 440
rect 229 -428 241 428
rect 275 -428 287 428
rect 229 -440 287 -428
rect 487 428 545 440
rect 487 -428 499 428
rect 533 -428 545 428
rect 487 -440 545 -428
rect 745 428 803 440
rect 745 -428 757 428
rect 791 -428 803 428
rect 745 -440 803 -428
rect 1003 428 1061 440
rect 1003 -428 1015 428
rect 1049 -428 1061 428
rect 1003 -440 1061 -428
rect 1261 428 1319 440
rect 1261 -428 1273 428
rect 1307 -428 1319 428
rect 1261 -440 1319 -428
rect 1519 428 1577 440
rect 1519 -428 1531 428
rect 1565 -428 1577 428
rect 1519 -440 1577 -428
rect 1777 428 1835 440
rect 1777 -428 1789 428
rect 1823 -428 1835 428
rect 1777 -440 1835 -428
<< mvndiffc >>
rect -1823 -428 -1789 428
rect -1565 -428 -1531 428
rect -1307 -428 -1273 428
rect -1049 -428 -1015 428
rect -791 -428 -757 428
rect -533 -428 -499 428
rect -275 -428 -241 428
rect -17 -428 17 428
rect 241 -428 275 428
rect 499 -428 533 428
rect 757 -428 791 428
rect 1015 -428 1049 428
rect 1273 -428 1307 428
rect 1531 -428 1565 428
rect 1789 -428 1823 428
<< mvpsubdiff >>
rect -1969 650 1969 662
rect -1969 616 -1861 650
rect 1861 616 1969 650
rect -1969 604 1969 616
rect -1969 554 -1911 604
rect -1969 -554 -1957 554
rect -1923 -554 -1911 554
rect 1911 554 1969 604
rect -1969 -604 -1911 -554
rect 1911 -554 1923 554
rect 1957 -554 1969 554
rect 1911 -604 1969 -554
rect -1969 -616 1969 -604
rect -1969 -650 -1861 -616
rect 1861 -650 1969 -616
rect -1969 -662 1969 -650
<< mvpsubdiffcont >>
rect -1861 616 1861 650
rect -1957 -554 -1923 554
rect 1923 -554 1957 554
rect -1861 -650 1861 -616
<< poly >>
rect -1777 512 -1577 528
rect -1777 478 -1761 512
rect -1593 478 -1577 512
rect -1777 440 -1577 478
rect -1519 512 -1319 528
rect -1519 478 -1503 512
rect -1335 478 -1319 512
rect -1519 440 -1319 478
rect -1261 512 -1061 528
rect -1261 478 -1245 512
rect -1077 478 -1061 512
rect -1261 440 -1061 478
rect -1003 512 -803 528
rect -1003 478 -987 512
rect -819 478 -803 512
rect -1003 440 -803 478
rect -745 512 -545 528
rect -745 478 -729 512
rect -561 478 -545 512
rect -745 440 -545 478
rect -487 512 -287 528
rect -487 478 -471 512
rect -303 478 -287 512
rect -487 440 -287 478
rect -229 512 -29 528
rect -229 478 -213 512
rect -45 478 -29 512
rect -229 440 -29 478
rect 29 512 229 528
rect 29 478 45 512
rect 213 478 229 512
rect 29 440 229 478
rect 287 512 487 528
rect 287 478 303 512
rect 471 478 487 512
rect 287 440 487 478
rect 545 512 745 528
rect 545 478 561 512
rect 729 478 745 512
rect 545 440 745 478
rect 803 512 1003 528
rect 803 478 819 512
rect 987 478 1003 512
rect 803 440 1003 478
rect 1061 512 1261 528
rect 1061 478 1077 512
rect 1245 478 1261 512
rect 1061 440 1261 478
rect 1319 512 1519 528
rect 1319 478 1335 512
rect 1503 478 1519 512
rect 1319 440 1519 478
rect 1577 512 1777 528
rect 1577 478 1593 512
rect 1761 478 1777 512
rect 1577 440 1777 478
rect -1777 -478 -1577 -440
rect -1777 -512 -1761 -478
rect -1593 -512 -1577 -478
rect -1777 -528 -1577 -512
rect -1519 -478 -1319 -440
rect -1519 -512 -1503 -478
rect -1335 -512 -1319 -478
rect -1519 -528 -1319 -512
rect -1261 -478 -1061 -440
rect -1261 -512 -1245 -478
rect -1077 -512 -1061 -478
rect -1261 -528 -1061 -512
rect -1003 -478 -803 -440
rect -1003 -512 -987 -478
rect -819 -512 -803 -478
rect -1003 -528 -803 -512
rect -745 -478 -545 -440
rect -745 -512 -729 -478
rect -561 -512 -545 -478
rect -745 -528 -545 -512
rect -487 -478 -287 -440
rect -487 -512 -471 -478
rect -303 -512 -287 -478
rect -487 -528 -287 -512
rect -229 -478 -29 -440
rect -229 -512 -213 -478
rect -45 -512 -29 -478
rect -229 -528 -29 -512
rect 29 -478 229 -440
rect 29 -512 45 -478
rect 213 -512 229 -478
rect 29 -528 229 -512
rect 287 -478 487 -440
rect 287 -512 303 -478
rect 471 -512 487 -478
rect 287 -528 487 -512
rect 545 -478 745 -440
rect 545 -512 561 -478
rect 729 -512 745 -478
rect 545 -528 745 -512
rect 803 -478 1003 -440
rect 803 -512 819 -478
rect 987 -512 1003 -478
rect 803 -528 1003 -512
rect 1061 -478 1261 -440
rect 1061 -512 1077 -478
rect 1245 -512 1261 -478
rect 1061 -528 1261 -512
rect 1319 -478 1519 -440
rect 1319 -512 1335 -478
rect 1503 -512 1519 -478
rect 1319 -528 1519 -512
rect 1577 -478 1777 -440
rect 1577 -512 1593 -478
rect 1761 -512 1777 -478
rect 1577 -528 1777 -512
<< polycont >>
rect -1761 478 -1593 512
rect -1503 478 -1335 512
rect -1245 478 -1077 512
rect -987 478 -819 512
rect -729 478 -561 512
rect -471 478 -303 512
rect -213 478 -45 512
rect 45 478 213 512
rect 303 478 471 512
rect 561 478 729 512
rect 819 478 987 512
rect 1077 478 1245 512
rect 1335 478 1503 512
rect 1593 478 1761 512
rect -1761 -512 -1593 -478
rect -1503 -512 -1335 -478
rect -1245 -512 -1077 -478
rect -987 -512 -819 -478
rect -729 -512 -561 -478
rect -471 -512 -303 -478
rect -213 -512 -45 -478
rect 45 -512 213 -478
rect 303 -512 471 -478
rect 561 -512 729 -478
rect 819 -512 987 -478
rect 1077 -512 1245 -478
rect 1335 -512 1503 -478
rect 1593 -512 1761 -478
<< locali >>
rect -1957 616 -1861 650
rect 1861 616 1957 650
rect -1957 554 -1923 616
rect 1923 554 1957 616
rect -1777 478 -1761 512
rect -1593 478 -1577 512
rect -1519 478 -1503 512
rect -1335 478 -1319 512
rect -1261 478 -1245 512
rect -1077 478 -1061 512
rect -1003 478 -987 512
rect -819 478 -803 512
rect -745 478 -729 512
rect -561 478 -545 512
rect -487 478 -471 512
rect -303 478 -287 512
rect -229 478 -213 512
rect -45 478 -29 512
rect 29 478 45 512
rect 213 478 229 512
rect 287 478 303 512
rect 471 478 487 512
rect 545 478 561 512
rect 729 478 745 512
rect 803 478 819 512
rect 987 478 1003 512
rect 1061 478 1077 512
rect 1245 478 1261 512
rect 1319 478 1335 512
rect 1503 478 1519 512
rect 1577 478 1593 512
rect 1761 478 1777 512
rect -1823 428 -1789 444
rect -1823 -444 -1789 -428
rect -1565 428 -1531 444
rect -1565 -444 -1531 -428
rect -1307 428 -1273 444
rect -1307 -444 -1273 -428
rect -1049 428 -1015 444
rect -1049 -444 -1015 -428
rect -791 428 -757 444
rect -791 -444 -757 -428
rect -533 428 -499 444
rect -533 -444 -499 -428
rect -275 428 -241 444
rect -275 -444 -241 -428
rect -17 428 17 444
rect -17 -444 17 -428
rect 241 428 275 444
rect 241 -444 275 -428
rect 499 428 533 444
rect 499 -444 533 -428
rect 757 428 791 444
rect 757 -444 791 -428
rect 1015 428 1049 444
rect 1015 -444 1049 -428
rect 1273 428 1307 444
rect 1273 -444 1307 -428
rect 1531 428 1565 444
rect 1531 -444 1565 -428
rect 1789 428 1823 444
rect 1789 -444 1823 -428
rect -1777 -512 -1761 -478
rect -1593 -512 -1577 -478
rect -1519 -512 -1503 -478
rect -1335 -512 -1319 -478
rect -1261 -512 -1245 -478
rect -1077 -512 -1061 -478
rect -1003 -512 -987 -478
rect -819 -512 -803 -478
rect -745 -512 -729 -478
rect -561 -512 -545 -478
rect -487 -512 -471 -478
rect -303 -512 -287 -478
rect -229 -512 -213 -478
rect -45 -512 -29 -478
rect 29 -512 45 -478
rect 213 -512 229 -478
rect 287 -512 303 -478
rect 471 -512 487 -478
rect 545 -512 561 -478
rect 729 -512 745 -478
rect 803 -512 819 -478
rect 987 -512 1003 -478
rect 1061 -512 1077 -478
rect 1245 -512 1261 -478
rect 1319 -512 1335 -478
rect 1503 -512 1519 -478
rect 1577 -512 1593 -478
rect 1761 -512 1777 -478
rect -1957 -616 -1923 -554
rect 1923 -616 1957 -554
rect -1957 -650 -1861 -616
rect 1861 -650 1957 -616
<< viali >>
rect -1761 478 -1593 512
rect -1503 478 -1335 512
rect -1245 478 -1077 512
rect -987 478 -819 512
rect -729 478 -561 512
rect -471 478 -303 512
rect -213 478 -45 512
rect 45 478 213 512
rect 303 478 471 512
rect 561 478 729 512
rect 819 478 987 512
rect 1077 478 1245 512
rect 1335 478 1503 512
rect 1593 478 1761 512
rect -1823 -428 -1789 428
rect -1565 -428 -1531 428
rect -1307 -428 -1273 428
rect -1049 -428 -1015 428
rect -791 -428 -757 428
rect -533 -428 -499 428
rect -275 -428 -241 428
rect -17 -428 17 428
rect 241 -428 275 428
rect 499 -428 533 428
rect 757 -428 791 428
rect 1015 -428 1049 428
rect 1273 -428 1307 428
rect 1531 -428 1565 428
rect 1789 -428 1823 428
rect -1761 -512 -1593 -478
rect -1503 -512 -1335 -478
rect -1245 -512 -1077 -478
rect -987 -512 -819 -478
rect -729 -512 -561 -478
rect -471 -512 -303 -478
rect -213 -512 -45 -478
rect 45 -512 213 -478
rect 303 -512 471 -478
rect 561 -512 729 -478
rect 819 -512 987 -478
rect 1077 -512 1245 -478
rect 1335 -512 1503 -478
rect 1593 -512 1761 -478
<< metal1 >>
rect -1773 512 -1581 518
rect -1773 478 -1761 512
rect -1593 478 -1581 512
rect -1773 472 -1581 478
rect -1515 512 -1323 518
rect -1515 478 -1503 512
rect -1335 478 -1323 512
rect -1515 472 -1323 478
rect -1257 512 -1065 518
rect -1257 478 -1245 512
rect -1077 478 -1065 512
rect -1257 472 -1065 478
rect -999 512 -807 518
rect -999 478 -987 512
rect -819 478 -807 512
rect -999 472 -807 478
rect -741 512 -549 518
rect -741 478 -729 512
rect -561 478 -549 512
rect -741 472 -549 478
rect -483 512 -291 518
rect -483 478 -471 512
rect -303 478 -291 512
rect -483 472 -291 478
rect -225 512 -33 518
rect -225 478 -213 512
rect -45 478 -33 512
rect -225 472 -33 478
rect 33 512 225 518
rect 33 478 45 512
rect 213 478 225 512
rect 33 472 225 478
rect 291 512 483 518
rect 291 478 303 512
rect 471 478 483 512
rect 291 472 483 478
rect 549 512 741 518
rect 549 478 561 512
rect 729 478 741 512
rect 549 472 741 478
rect 807 512 999 518
rect 807 478 819 512
rect 987 478 999 512
rect 807 472 999 478
rect 1065 512 1257 518
rect 1065 478 1077 512
rect 1245 478 1257 512
rect 1065 472 1257 478
rect 1323 512 1515 518
rect 1323 478 1335 512
rect 1503 478 1515 512
rect 1323 472 1515 478
rect 1581 512 1773 518
rect 1581 478 1593 512
rect 1761 478 1773 512
rect 1581 472 1773 478
rect -1829 428 -1783 440
rect -1829 -428 -1823 428
rect -1789 -428 -1783 428
rect -1829 -440 -1783 -428
rect -1571 428 -1525 440
rect -1571 -428 -1565 428
rect -1531 -428 -1525 428
rect -1571 -440 -1525 -428
rect -1313 428 -1267 440
rect -1313 -428 -1307 428
rect -1273 -428 -1267 428
rect -1313 -440 -1267 -428
rect -1055 428 -1009 440
rect -1055 -428 -1049 428
rect -1015 -428 -1009 428
rect -1055 -440 -1009 -428
rect -797 428 -751 440
rect -797 -428 -791 428
rect -757 -428 -751 428
rect -797 -440 -751 -428
rect -539 428 -493 440
rect -539 -428 -533 428
rect -499 -428 -493 428
rect -539 -440 -493 -428
rect -281 428 -235 440
rect -281 -428 -275 428
rect -241 -428 -235 428
rect -281 -440 -235 -428
rect -23 428 23 440
rect -23 -428 -17 428
rect 17 -428 23 428
rect -23 -440 23 -428
rect 235 428 281 440
rect 235 -428 241 428
rect 275 -428 281 428
rect 235 -440 281 -428
rect 493 428 539 440
rect 493 -428 499 428
rect 533 -428 539 428
rect 493 -440 539 -428
rect 751 428 797 440
rect 751 -428 757 428
rect 791 -428 797 428
rect 751 -440 797 -428
rect 1009 428 1055 440
rect 1009 -428 1015 428
rect 1049 -428 1055 428
rect 1009 -440 1055 -428
rect 1267 428 1313 440
rect 1267 -428 1273 428
rect 1307 -428 1313 428
rect 1267 -440 1313 -428
rect 1525 428 1571 440
rect 1525 -428 1531 428
rect 1565 -428 1571 428
rect 1525 -440 1571 -428
rect 1783 428 1829 440
rect 1783 -428 1789 428
rect 1823 -428 1829 428
rect 1783 -440 1829 -428
rect -1773 -478 -1581 -472
rect -1773 -512 -1761 -478
rect -1593 -512 -1581 -478
rect -1773 -518 -1581 -512
rect -1515 -478 -1323 -472
rect -1515 -512 -1503 -478
rect -1335 -512 -1323 -478
rect -1515 -518 -1323 -512
rect -1257 -478 -1065 -472
rect -1257 -512 -1245 -478
rect -1077 -512 -1065 -478
rect -1257 -518 -1065 -512
rect -999 -478 -807 -472
rect -999 -512 -987 -478
rect -819 -512 -807 -478
rect -999 -518 -807 -512
rect -741 -478 -549 -472
rect -741 -512 -729 -478
rect -561 -512 -549 -478
rect -741 -518 -549 -512
rect -483 -478 -291 -472
rect -483 -512 -471 -478
rect -303 -512 -291 -478
rect -483 -518 -291 -512
rect -225 -478 -33 -472
rect -225 -512 -213 -478
rect -45 -512 -33 -478
rect -225 -518 -33 -512
rect 33 -478 225 -472
rect 33 -512 45 -478
rect 213 -512 225 -478
rect 33 -518 225 -512
rect 291 -478 483 -472
rect 291 -512 303 -478
rect 471 -512 483 -478
rect 291 -518 483 -512
rect 549 -478 741 -472
rect 549 -512 561 -478
rect 729 -512 741 -478
rect 549 -518 741 -512
rect 807 -478 999 -472
rect 807 -512 819 -478
rect 987 -512 999 -478
rect 807 -518 999 -512
rect 1065 -478 1257 -472
rect 1065 -512 1077 -478
rect 1245 -512 1257 -478
rect 1065 -518 1257 -512
rect 1323 -478 1515 -472
rect 1323 -512 1335 -478
rect 1503 -512 1515 -478
rect 1323 -518 1515 -512
rect 1581 -478 1773 -472
rect 1581 -512 1593 -478
rect 1761 -512 1773 -478
rect 1581 -518 1773 -512
<< properties >>
string FIXED_BBOX -1940 -633 1940 633
string gencell sky130_fd_pr__nfet_g5v0d10v5
string library sky130
string parameters w 4.4 l 1.0 m 1 nf 14 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
