magic
tech sky130A
timestamp 1716973465
<< end >>
