** sch_path: /home/tim/gits/cheetah_v3_analog/dependencies/sky130_hcmus_ip__instramp/cace/templates/dccurrent_vdd.sch
**.subckt dccurrent_vdd
VVcm net3 VSUB DC {Vcm}
Vena ena VSUB DC [{ena} * {Vdvdd}]
Vvss vss VSUB DC {Vvss}
Rout out VSUB {Rout} m=1
Cout out VSUB {Cout} m=1
Vvdd vdd VSUB DC {Vvdd}
RSUB VSUB GND 0.01 m=1
VVdiff net3 inp DC [{Vdiff} / 2]
x2 vdd vss net3 inm inp d0 d1 d2 d3 d4 d5 d6 d7 d8 d9 net2 net1 out ibias ena DVDD vss sky130_hcmus_ip__instramp
* noconn #net2
* noconn #net1
VDVDD1 DVDD VSUB DC {Vdvdd}
Iibias VSUB ibias {Ibias}
Vd0 d0 VSUB DC [{D[0]} * {Vdvdd}]
Vd1 d1 VSUB DC [{D[1]} * {Vdvdd}]
Vd2 d2 VSUB DC [{D[2]} * {Vdvdd}]
Vd3 d3 VSUB DC [{D[3]} * {Vdvdd}]
Vd4 d4 VSUB DC [{D[4]} * {Vdvdd}]
Vd5 d5 VSUB DC [{D[5]} * {Vdvdd}]
Vd6 d6 VSUB DC [{D[6]} * {Vdvdd}]
Vd7 d7 VSUB DC [{D[7]} * {Vdvdd}]
Vd8 d8 VSUB DC [{D[8]} * {Vdvdd}]
Vd9 d9 VSUB DC [{D[9]} * {Vdvdd}]
VVdiff1 inm net3 DC [{Vdiff} / 2]
**** begin user architecture code

.control
op
set wr_singlescale
wrdata {simpath}/{filename}_{N}.data -I(Vvdd)
quit
.endc



* CACE gensim simulation file {filename}_{N}
* Generated by CACE gensim, Efabless Corporation (c) 2023
* Find the noise in the driver amplifier

.include {DUT_path}

.lib {PDK_ROOT}/{PDK}/libs.tech/combined/sky130.lib.spice {corner}
.include {PDK_ROOT}/{PDK}/libs.ref/sky130_fd_sc_hvl/spice/sky130_fd_sc_hvl.spice

.option TEMP={temperature}
* Flag unsafe operating conditions (exceeds models' specified limits)
.option warn=1


**** end user architecture code
**.ends
.GLOBAL GND
.end
