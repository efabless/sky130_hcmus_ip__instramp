* NGSPICE file created from sky130_hcmus_ip__instramp.ext - technology: sky130A

.subckt sky130_fd_pr__res_high_po_0p69_JKKHRG a_n199_n1768# a_n69_1206# a_n69_n1638#
X0 a_n69_1206# a_n69_n1638# a_n199_n1768# sky130_fd_pr__res_high_po_0p69 l=12.22
.ends

.subckt sky130_fd_pr__res_high_po_0p69_Z3RMRJ a_48_1206# a_n186_n1638# a_n186_1206#
+ a_n316_n1768# a_48_n1638#
X0 a_48_1206# a_48_n1638# a_n316_n1768# sky130_fd_pr__res_high_po_0p69 l=12.22
X1 a_n186_1206# a_n186_n1638# a_n316_n1768# sky130_fd_pr__res_high_po_0p69 l=12.22
.ends

.subckt sky130_fd_pr__res_high_po_0p69_Z3RMR6 a_516_n1638# a_48_1206# a_n654_1206#
+ a_n888_1206# a_n186_n1638# a_n186_1206# a_750_1206# a_n654_n1638# a_282_1206# a_282_n1638#
+ a_48_n1638# a_750_n1638# a_n420_n1638# a_516_1206# a_n1018_n1768# a_n420_1206# a_n888_n1638#
X0 a_n420_1206# a_n420_n1638# a_n1018_n1768# sky130_fd_pr__res_high_po_0p69 l=12.22
X1 a_48_1206# a_48_n1638# a_n1018_n1768# sky130_fd_pr__res_high_po_0p69 l=12.22
X2 a_750_1206# a_750_n1638# a_n1018_n1768# sky130_fd_pr__res_high_po_0p69 l=12.22
X3 a_n888_1206# a_n888_n1638# a_n1018_n1768# sky130_fd_pr__res_high_po_0p69 l=12.22
X4 a_282_1206# a_282_n1638# a_n1018_n1768# sky130_fd_pr__res_high_po_0p69 l=12.22
X5 a_n654_1206# a_n654_n1638# a_n1018_n1768# sky130_fd_pr__res_high_po_0p69 l=12.22
X6 a_n186_1206# a_n186_n1638# a_n1018_n1768# sky130_fd_pr__res_high_po_0p69 l=12.22
X7 a_516_1206# a_516_n1638# a_n1018_n1768# sky130_fd_pr__res_high_po_0p69 l=12.22
.ends

.subckt sky130_fd_pr__res_high_po_0p69_YMHKRJ a_48_1206# a_n550_n1768# a_n186_n1638#
+ a_n186_1206# a_282_1206# a_282_n1638# a_48_n1638# a_n420_n1638# a_n420_1206#
X0 a_n420_1206# a_n420_n1638# a_n550_n1768# sky130_fd_pr__res_high_po_0p69 l=12.22
X1 a_48_1206# a_48_n1638# a_n550_n1768# sky130_fd_pr__res_high_po_0p69 l=12.22
X2 a_282_1206# a_282_n1638# a_n550_n1768# sky130_fd_pr__res_high_po_0p69 l=12.22
X3 a_n186_1206# a_n186_n1638# a_n550_n1768# sky130_fd_pr__res_high_po_0p69 l=12.22
.ends

.subckt sky130_fd_pr__res_high_po_0p69_HBQF5Z a_516_n1638# a_48_1206# a_n654_1206#
+ a_n888_1206# a_1452_1206# a_n1122_n1638# a_1452_n1638# a_n186_n1638# a_n186_1206#
+ a_n1954_n1768# a_1686_1206# a_750_1206# a_n654_n1638# a_n1590_1206# a_984_n1638#
+ a_984_1206# a_n1824_1206# a_n1590_n1638# a_1218_n1638# a_282_1206# a_n1122_1206#
+ a_1218_1206# a_282_n1638# a_48_n1638# a_750_n1638# a_n420_n1638# a_n1356_1206# a_516_1206#
+ a_n1356_n1638# a_1686_n1638# a_n420_1206# a_n1824_n1638# a_n888_n1638#
X0 a_n420_1206# a_n420_n1638# a_n1954_n1768# sky130_fd_pr__res_high_po_0p69 l=12.22
X1 a_1452_1206# a_1452_n1638# a_n1954_n1768# sky130_fd_pr__res_high_po_0p69 l=12.22
X2 a_n1824_1206# a_n1824_n1638# a_n1954_n1768# sky130_fd_pr__res_high_po_0p69 l=12.22
X3 a_n1590_1206# a_n1590_n1638# a_n1954_n1768# sky130_fd_pr__res_high_po_0p69 l=12.22
X4 a_48_1206# a_48_n1638# a_n1954_n1768# sky130_fd_pr__res_high_po_0p69 l=12.22
X5 a_984_1206# a_984_n1638# a_n1954_n1768# sky130_fd_pr__res_high_po_0p69 l=12.22
X6 a_n1356_1206# a_n1356_n1638# a_n1954_n1768# sky130_fd_pr__res_high_po_0p69 l=12.22
X7 a_1218_1206# a_1218_n1638# a_n1954_n1768# sky130_fd_pr__res_high_po_0p69 l=12.22
X8 a_750_1206# a_750_n1638# a_n1954_n1768# sky130_fd_pr__res_high_po_0p69 l=12.22
X9 a_n1122_1206# a_n1122_n1638# a_n1954_n1768# sky130_fd_pr__res_high_po_0p69 l=12.22
X10 a_n888_1206# a_n888_n1638# a_n1954_n1768# sky130_fd_pr__res_high_po_0p69 l=12.22
X11 a_282_1206# a_282_n1638# a_n1954_n1768# sky130_fd_pr__res_high_po_0p69 l=12.22
X12 a_n654_1206# a_n654_n1638# a_n1954_n1768# sky130_fd_pr__res_high_po_0p69 l=12.22
X13 a_n186_1206# a_n186_n1638# a_n1954_n1768# sky130_fd_pr__res_high_po_0p69 l=12.22
X14 a_516_1206# a_516_n1638# a_n1954_n1768# sky130_fd_pr__res_high_po_0p69 l=12.22
X15 a_1686_1206# a_1686_n1638# a_n1954_n1768# sky130_fd_pr__res_high_po_0p69 l=12.22
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_727CUP a_n100_n565# a_100_n477# a_n292_n699#
+ a_n158_n477#
X0 a_100_n477# a_n100_n565# a_n158_n477# a_n292_n699# sky130_fd_pr__nfet_g5v0d10v5 ad=1.3833 pd=10.12 as=1.3833 ps=10.12 w=4.77 l=1
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_VU5C5A a_n287_n487# a_n421_n709# a_n229_n575#
+ a_229_n487# a_n29_n487# a_29_n575#
X0 a_229_n487# a_29_n575# a_n29_n487# a_n421_n709# sky130_fd_pr__nfet_g5v0d10v5 ad=1.4123 pd=10.32 as=0.70615 ps=5.16 w=4.87 l=1
X1 a_n29_n487# a_n229_n575# a_n287_n487# a_n421_n709# sky130_fd_pr__nfet_g5v0d10v5 ad=0.70615 pd=5.16 as=1.4123 ps=10.32 w=4.87 l=1
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_J97EKB a_487_n438# a_n803_n438# a_29_n526# a_n745_n526#
+ a_n287_n438# a_n1061_n438# a_803_n526# a_745_n438# a_n229_n526# a_287_n526# a_n1003_n526#
+ a_229_n438# a_n545_n438# a_1003_n438# a_n487_n526# a_n1195_n660# a_545_n526# a_n29_n438#
X0 a_1003_n438# a_803_n526# a_745_n438# a_n1195_n660# sky130_fd_pr__nfet_g5v0d10v5 ad=1.2702 pd=9.34 as=0.6351 ps=4.67 w=4.38 l=1
X1 a_745_n438# a_545_n526# a_487_n438# a_n1195_n660# sky130_fd_pr__nfet_g5v0d10v5 ad=0.6351 pd=4.67 as=0.6351 ps=4.67 w=4.38 l=1
X2 a_487_n438# a_287_n526# a_229_n438# a_n1195_n660# sky130_fd_pr__nfet_g5v0d10v5 ad=0.6351 pd=4.67 as=0.6351 ps=4.67 w=4.38 l=1
X3 a_229_n438# a_29_n526# a_n29_n438# a_n1195_n660# sky130_fd_pr__nfet_g5v0d10v5 ad=0.6351 pd=4.67 as=0.6351 ps=4.67 w=4.38 l=1
X4 a_n29_n438# a_n229_n526# a_n287_n438# a_n1195_n660# sky130_fd_pr__nfet_g5v0d10v5 ad=0.6351 pd=4.67 as=0.6351 ps=4.67 w=4.38 l=1
X5 a_n545_n438# a_n745_n526# a_n803_n438# a_n1195_n660# sky130_fd_pr__nfet_g5v0d10v5 ad=0.6351 pd=4.67 as=0.6351 ps=4.67 w=4.38 l=1
X6 a_n287_n438# a_n487_n526# a_n545_n438# a_n1195_n660# sky130_fd_pr__nfet_g5v0d10v5 ad=0.6351 pd=4.67 as=0.6351 ps=4.67 w=4.38 l=1
X7 a_n803_n438# a_n1003_n526# a_n1061_n438# a_n1195_n660# sky130_fd_pr__nfet_g5v0d10v5 ad=0.6351 pd=4.67 as=1.2702 ps=9.34 w=4.38 l=1
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_S7E57E a_n229_n553# a_287_n553# a_229_n465# a_n545_n465#
+ a_n487_n553# a_487_n465# a_n29_n465# a_n679_n687# a_29_n553# a_n287_n465#
X0 a_487_n465# a_287_n553# a_229_n465# a_n679_n687# sky130_fd_pr__nfet_g5v0d10v5 ad=1.3485 pd=9.88 as=0.67425 ps=4.94 w=4.65 l=1
X1 a_229_n465# a_29_n553# a_n29_n465# a_n679_n687# sky130_fd_pr__nfet_g5v0d10v5 ad=0.67425 pd=4.94 as=0.67425 ps=4.94 w=4.65 l=1
X2 a_n29_n465# a_n229_n553# a_n287_n465# a_n679_n687# sky130_fd_pr__nfet_g5v0d10v5 ad=0.67425 pd=4.94 as=0.67425 ps=4.94 w=4.65 l=1
X3 a_n287_n465# a_n487_n553# a_n545_n465# a_n679_n687# sky130_fd_pr__nfet_g5v0d10v5 ad=0.67425 pd=4.94 as=1.3485 ps=9.88 w=4.65 l=1
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_YPGNM4 a_545_n528# a_n545_n440# a_1577_n528#
+ a_1003_n440# a_n29_n440# a_29_n528# a_n1777_n528# a_487_n440# a_n745_n528# a_n1835_n440#
+ a_803_n528# a_n803_n440# a_1519_n440# a_1261_n440# a_n229_n528# a_n1319_n440# a_287_n528#
+ a_n1003_n528# a_n287_n440# a_n1061_n440# a_n1969_n662# a_745_n440# a_1319_n528#
+ a_1061_n528# a_1777_n440# a_n1519_n528# a_229_n440# a_n487_n528# a_n1261_n528# a_n1577_n440#
X0 a_1777_n440# a_1577_n528# a_1519_n440# a_n1969_n662# sky130_fd_pr__nfet_g5v0d10v5 ad=1.276 pd=9.38 as=0.638 ps=4.69 w=4.4 l=1
X1 a_1261_n440# a_1061_n528# a_1003_n440# a_n1969_n662# sky130_fd_pr__nfet_g5v0d10v5 ad=0.638 pd=4.69 as=0.638 ps=4.69 w=4.4 l=1
X2 a_229_n440# a_29_n528# a_n29_n440# a_n1969_n662# sky130_fd_pr__nfet_g5v0d10v5 ad=0.638 pd=4.69 as=0.638 ps=4.69 w=4.4 l=1
X3 a_n29_n440# a_n229_n528# a_n287_n440# a_n1969_n662# sky130_fd_pr__nfet_g5v0d10v5 ad=0.638 pd=4.69 as=0.638 ps=4.69 w=4.4 l=1
X4 a_n1319_n440# a_n1519_n528# a_n1577_n440# a_n1969_n662# sky130_fd_pr__nfet_g5v0d10v5 ad=0.638 pd=4.69 as=0.638 ps=4.69 w=4.4 l=1
X5 a_n545_n440# a_n745_n528# a_n803_n440# a_n1969_n662# sky130_fd_pr__nfet_g5v0d10v5 ad=0.638 pd=4.69 as=0.638 ps=4.69 w=4.4 l=1
X6 a_n803_n440# a_n1003_n528# a_n1061_n440# a_n1969_n662# sky130_fd_pr__nfet_g5v0d10v5 ad=0.638 pd=4.69 as=0.638 ps=4.69 w=4.4 l=1
X7 a_n287_n440# a_n487_n528# a_n545_n440# a_n1969_n662# sky130_fd_pr__nfet_g5v0d10v5 ad=0.638 pd=4.69 as=0.638 ps=4.69 w=4.4 l=1
X8 a_n1577_n440# a_n1777_n528# a_n1835_n440# a_n1969_n662# sky130_fd_pr__nfet_g5v0d10v5 ad=0.638 pd=4.69 as=1.276 ps=9.38 w=4.4 l=1
X9 a_1519_n440# a_1319_n528# a_1261_n440# a_n1969_n662# sky130_fd_pr__nfet_g5v0d10v5 ad=0.638 pd=4.69 as=0.638 ps=4.69 w=4.4 l=1
X10 a_n1061_n440# a_n1261_n528# a_n1319_n440# a_n1969_n662# sky130_fd_pr__nfet_g5v0d10v5 ad=0.638 pd=4.69 as=0.638 ps=4.69 w=4.4 l=1
X11 a_1003_n440# a_803_n528# a_745_n440# a_n1969_n662# sky130_fd_pr__nfet_g5v0d10v5 ad=0.638 pd=4.69 as=0.638 ps=4.69 w=4.4 l=1
X12 a_487_n440# a_287_n528# a_229_n440# a_n1969_n662# sky130_fd_pr__nfet_g5v0d10v5 ad=0.638 pd=4.69 as=0.638 ps=4.69 w=4.4 l=1
X13 a_745_n440# a_545_n528# a_487_n440# a_n1969_n662# sky130_fd_pr__nfet_g5v0d10v5 ad=0.638 pd=4.69 as=0.638 ps=4.69 w=4.4 l=1
.ends

.subckt RB_array_20 VDD R1 D0 D3 D4 R2 D1 D2 VSS
XXR1 VSS R2 m1_2651_1472# sky130_fd_pr__res_high_po_0p69_JKKHRG
XXR2 VSS R2 m1_2124_1470# sky130_fd_pr__res_high_po_0p69_JKKHRG
XXR3 R2 m1_3160_410# R2 VSS m1_3160_410# sky130_fd_pr__res_high_po_0p69_Z3RMRJ
XXR5 m1_5470_410# R2 R2 R2 m1_5470_410# R2 R2 m1_5470_410# R2 m1_5470_410# m1_5470_410#
+ m1_5470_410# m1_5470_410# R2 VSS R2 m1_5470_410# sky130_fd_pr__res_high_po_0p69_Z3RMR6
XXR4 R2 VSS m1_4060_410# R2 R2 m1_4060_410# m1_4060_410# m1_4060_410# R2 sky130_fd_pr__res_high_po_0p69_YMHKRJ
XXR6 m1_7940_410# R2 R2 R2 R2 m1_7940_410# m1_7940_410# m1_7940_410# R2 VSS R2 R2
+ m1_7940_410# R2 m1_7940_410# R2 R2 m1_7940_410# m1_7940_410# R2 R2 R2 m1_7940_410#
+ m1_7940_410# m1_7940_410# m1_7940_410# R2 R2 m1_7940_410# m1_7940_410# R2 m1_7940_410#
+ m1_7940_410# sky130_fd_pr__res_high_po_0p69_HBQF5Z
XXM6 D0 m1_2651_1472# VSS R1 sky130_fd_pr__nfet_g5v0d10v5_727CUP
XXM7 m1_3160_410# VSS D1 m1_3160_410# R1 D1 sky130_fd_pr__nfet_g5v0d10v5_VU5C5A
XXM9 m1_5470_410# R1 D3 D3 R1 m1_5470_410# D3 R1 D3 D3 D3 R1 m1_5470_410# m1_5470_410#
+ D3 VSS D3 m1_5470_410# sky130_fd_pr__nfet_g5v0d10v5_J97EKB
XXM8 D2 D2 R1 m1_4060_410# D2 m1_4060_410# m1_4060_410# VSS D2 R1 sky130_fd_pr__nfet_g5v0d10v5_S7E57E
XXM10 D4 R1 D4 R1 R1 D4 D4 R1 D4 m1_7940_410# D4 m1_7940_410# R1 m1_7940_410# D4 m1_7940_410#
+ D4 D4 m1_7940_410# R1 VSS m1_7940_410# D4 D4 m1_7940_410# D4 m1_7940_410# D4 D4
+ R1 sky130_fd_pr__nfet_g5v0d10v5_YPGNM4
XXM11 VDD m1_2124_1470# VSS R1 sky130_fd_pr__nfet_g5v0d10v5_727CUP
.ends

.subckt sky130_fd_pr__res_high_po_0p69_T8KQH6 a_n199_n866# a_n69_n736# a_n69_304#
X0 a_n69_304# a_n69_n736# a_n199_n866# sky130_fd_pr__res_high_po_0p69 l=3.2
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_K8DQNF a_n29_n1536# a_229_n1536# a_n229_n1562#
+ w_n487_n1762# a_n287_n1536# a_29_n1562#
X0 a_n29_n1536# a_n229_n1562# a_n287_n1536# w_n487_n1762# sky130_fd_pr__pfet_g5v0d10v5 ad=2.175 pd=15.29 as=4.35 ps=30.58 w=15 l=1
X1 a_229_n1536# a_29_n1562# a_n29_n1536# w_n487_n1762# sky130_fd_pr__pfet_g5v0d10v5 ad=4.35 pd=30.58 as=2.175 ps=15.29 w=15 l=1
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_VYCZE8 a_100_n1681# a_n292_n1841# a_n100_n1707#
+ a_n158_n1681#
X0 a_100_n1681# a_n100_n1707# a_n158_n1681# a_n292_n1841# sky130_fd_pr__nfet_g5v0d10v5 ad=4.785 pd=33.58 as=4.785 ps=33.58 w=16.5 l=1
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_F3SB2X a_n100_n1632# a_100_n1544# a_n292_n1766#
+ a_n158_n1544#
X0 a_100_n1544# a_n100_n1632# a_n158_n1544# a_n292_n1766# sky130_fd_pr__nfet_g5v0d10v5 ad=4.4776 pd=31.46 as=4.4776 ps=31.46 w=15.44 l=1
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_2HXNYY a_n158_n1900# a_100_n1900# a_n292_n2122#
+ a_n100_n1988#
X0 a_100_n1900# a_n100_n1988# a_n158_n1900# a_n292_n2122# sky130_fd_pr__nfet_g5v0d10v5 ad=5.51 pd=38.58 as=5.51 ps=38.58 w=19 l=1
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_24QKAW a_29_n1997# a_n487_n1997# a_487_n1900#
+ a_n287_n1900# a_n229_n1997# a_n545_n1900# a_n29_n1900# a_287_n1997# w_n745_n2197#
+ a_229_n1900#
X0 a_487_n1900# a_287_n1997# a_229_n1900# w_n745_n2197# sky130_fd_pr__pfet_g5v0d10v5 ad=5.51 pd=38.58 as=2.755 ps=19.29 w=19 l=1
X1 a_n287_n1900# a_n487_n1997# a_n545_n1900# w_n745_n2197# sky130_fd_pr__pfet_g5v0d10v5 ad=2.755 pd=19.29 as=5.51 ps=38.58 w=19 l=1
X2 a_n29_n1900# a_n229_n1997# a_n287_n1900# w_n745_n2197# sky130_fd_pr__pfet_g5v0d10v5 ad=2.755 pd=19.29 as=2.755 ps=19.29 w=19 l=1
X3 a_229_n1900# a_29_n1997# a_n29_n1900# w_n745_n2197# sky130_fd_pr__pfet_g5v0d10v5 ad=2.755 pd=19.29 as=2.755 ps=19.29 w=19 l=1
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_LB7Y8R a_n100_n157# a_n158_n69# a_n292_n291#
+ a_100_n69#
X0 a_100_n69# a_n100_n157# a_n158_n69# a_n292_n291# sky130_fd_pr__nfet_g5v0d10v5 ad=0.2001 pd=1.96 as=0.2001 ps=1.96 w=0.69 l=1
.ends

.subckt sky130_fd_pr__cap_mim_m3_1_8DB3RK m3_n876_n730# c1_n836_n690#
X0 c1_n836_n690# m3_n876_n730# sky130_fd_pr__cap_mim_m3_1 l=6.9 w=6.9
.ends

.subckt opamp V1 V2 VOUT VDD VSS
XXR3 VSS m1_4128_540# VOUT sky130_fd_pr__res_high_po_0p69_T8KQH6
XXM1 m1_5053_7611# VDD a_4864_8007# VDD VDD a_4864_8007# sky130_fd_pr__pfet_g5v0d10v5_K8DQNF
XXM2 m1_4306_994# VSS V2 a_4864_8007# sky130_fd_pr__nfet_g5v0d10v5_VYCZE8
XXM3 a_4864_8007# VDD a_4864_8007# VDD VDD a_4864_8007# sky130_fd_pr__pfet_g5v0d10v5_K8DQNF
XXM4 m1_5053_7611# VSS V1 m1_4306_994# sky130_fd_pr__nfet_g5v0d10v5_VYCZE8
XXM5 m1_5284_1188# VSS VSS m1_4306_994# sky130_fd_pr__nfet_g5v0d10v5_F3SB2X
XXM6 VSS VOUT VSS m1_5284_1188# sky130_fd_pr__nfet_g5v0d10v5_2HXNYY
XXM7 m1_5284_1188# m1_5284_1188# VSS VSS sky130_fd_pr__nfet_g5v0d10v5_F3SB2X
XXM8 m1_5053_7611# m1_5053_7611# VDD VOUT m1_5053_7611# VDD VDD m1_5053_7611# VDD
+ VOUT sky130_fd_pr__pfet_g5v0d10v5_24QKAW
XXM9 VDD VDD VSS m1_5284_1188# sky130_fd_pr__nfet_g5v0d10v5_LB7Y8R
XXC1 m1_5053_7611# m1_4128_540# sky130_fd_pr__cap_mim_m3_1_8DB3RK
.ends

.subckt sky130_fd_pr__res_high_po_0p69_WX3C5M a_2856_n1638# a_3090_1206# a_n3930_1206#
+ a_n5100_n1638# a_4260_n1638# a_7068_1206# a_516_n1638# a_6600_1206# a_n654_1206#
+ a_48_1206# a_4728_n1638# a_5196_1206# a_6132_n1638# a_n2526_1206# a_n6972_n1638#
+ a_5430_n1638# a_n5100_1206# a_3324_1206# a_6834_1206# a_7302_n1638# a_6600_n1638#
+ a_n888_1206# a_n7206_1206# a_n1122_n1638# a_1452_1206# a_4962_1206# a_n5334_1206#
+ a_n4398_n1638# a_n186_n1638# a_n3696_n1638# a_n2994_n1638# a_2154_n1638# a_n3462_1206#
+ a_n6972_1206# a_1452_n1638# a_3558_1206# a_6132_1206# a_n186_1206# a_n5568_n1638#
+ a_n1590_1206# a_n4866_n1638# a_1686_1206# a_4026_n1638# a_750_1206# a_3324_n1638#
+ a_n654_n1638# a_n2058_1206# a_n5568_1206# a_n6270_n1638# a_4260_1206# a_2622_n1638#
+ a_1920_n1638# a_984_n1638# a_n6738_n1638# a_n3696_1206# a_5898_n1638# a_n6270_1206#
+ a_6366_1206# a_n7440_n1638# a_984_1206# a_4494_1206# a_n1824_1206# a_n2292_n1638#
+ a_n1590_n1638# a_2622_1206# a_n6504_1206# a_1218_n1638# a_282_1206# a_n4164_n1638#
+ a_n3462_n1638# a_n2760_n1638# a_n1122_1206# a_n4632_1206# a_282_n1638# a_1218_1206#
+ a_4728_1206# a_7302_1206# a_n6036_n1638# a_5196_n1638# a_n5334_n1638# a_48_n1638#
+ a_n2760_1206# a_2856_1206# a_4494_n1638# a_n4632_n1638# a_3792_n1638# a_n3228_1206#
+ a_n3930_n1638# a_n6738_1206# a_n420_n1638# a_5430_1206# a_750_n1638# a_7068_n1638#
+ a_n7206_n1638# a_6366_n1638# a_n1356_1206# a_n4866_1206# a_n6504_n1638# a_5664_n1638#
+ a_n5802_n1638# a_516_1206# a_n7440_1206# a_4962_n1638# a_4026_1206# a_n7570_n1768#
+ a_n2994_1206# a_2154_1206# a_5664_1206# a_6834_n1638# a_n6036_1206# a_n2058_n1638#
+ a_n1356_n1638# a_3792_1206# a_n4164_1206# a_n3228_n1638# a_2388_n1638# a_n2526_n1638#
+ a_n420_1206# a_n2292_1206# a_1686_n1638# a_2388_1206# a_5898_1206# a_n1824_n1638#
+ a_3090_n1638# a_1920_1206# a_n5802_1206# a_3558_n1638# a_n888_n1638# a_n4398_1206#
X0 a_n420_1206# a_n420_n1638# a_n7570_n1768# sky130_fd_pr__res_high_po_0p69 l=12.22
X1 a_3090_1206# a_3090_n1638# a_n7570_n1768# sky130_fd_pr__res_high_po_0p69 l=12.22
X2 a_n6036_1206# a_n6036_n1638# a_n7570_n1768# sky130_fd_pr__res_high_po_0p69 l=12.22
X3 a_n2058_1206# a_n2058_n1638# a_n7570_n1768# sky130_fd_pr__res_high_po_0p69 l=12.22
X4 a_1452_1206# a_1452_n1638# a_n7570_n1768# sky130_fd_pr__res_high_po_0p69 l=12.22
X5 a_5430_1206# a_5430_n1638# a_n7570_n1768# sky130_fd_pr__res_high_po_0p69 l=12.22
X6 a_5196_1206# a_5196_n1638# a_n7570_n1768# sky130_fd_pr__res_high_po_0p69 l=12.22
X7 a_n3696_1206# a_n3696_n1638# a_n7570_n1768# sky130_fd_pr__res_high_po_0p69 l=12.22
X8 a_3558_1206# a_3558_n1638# a_n7570_n1768# sky130_fd_pr__res_high_po_0p69 l=12.22
X9 a_n3462_1206# a_n3462_n1638# a_n7570_n1768# sky130_fd_pr__res_high_po_0p69 l=12.22
X10 a_3324_1206# a_3324_n1638# a_n7570_n1768# sky130_fd_pr__res_high_po_0p69 l=12.22
X11 a_7068_1206# a_7068_n1638# a_n7570_n1768# sky130_fd_pr__res_high_po_0p69 l=12.22
X12 a_7302_1206# a_7302_n1638# a_n7570_n1768# sky130_fd_pr__res_high_po_0p69 l=12.22
X13 a_n5802_1206# a_n5802_n1638# a_n7570_n1768# sky130_fd_pr__res_high_po_0p69 l=12.22
X14 a_n1824_1206# a_n1824_n1638# a_n7570_n1768# sky130_fd_pr__res_high_po_0p69 l=12.22
X15 a_n5568_1206# a_n5568_n1638# a_n7570_n1768# sky130_fd_pr__res_high_po_0p69 l=12.22
X16 a_n1590_1206# a_n1590_n1638# a_n7570_n1768# sky130_fd_pr__res_high_po_0p69 l=12.22
X17 a_4962_1206# a_4962_n1638# a_n7570_n1768# sky130_fd_pr__res_high_po_0p69 l=12.22
X18 a_48_1206# a_48_n1638# a_n7570_n1768# sky130_fd_pr__res_high_po_0p69 l=12.22
X19 a_n3930_1206# a_n3930_n1638# a_n7570_n1768# sky130_fd_pr__res_high_po_0p69 l=12.22
X20 a_984_1206# a_984_n1638# a_n7570_n1768# sky130_fd_pr__res_high_po_0p69 l=12.22
X21 a_n5334_1206# a_n5334_n1638# a_n7570_n1768# sky130_fd_pr__res_high_po_0p69 l=12.22
X22 a_n1356_1206# a_n1356_n1638# a_n7570_n1768# sky130_fd_pr__res_high_po_0p69 l=12.22
X23 a_n5100_1206# a_n5100_n1638# a_n7570_n1768# sky130_fd_pr__res_high_po_0p69 l=12.22
X24 a_1218_1206# a_1218_n1638# a_n7570_n1768# sky130_fd_pr__res_high_po_0p69 l=12.22
X25 a_4494_1206# a_4494_n1638# a_n7570_n1768# sky130_fd_pr__res_high_po_0p69 l=12.22
X26 a_n6972_1206# a_n6972_n1638# a_n7570_n1768# sky130_fd_pr__res_high_po_0p69 l=12.22
X27 a_n2994_1206# a_n2994_n1638# a_n7570_n1768# sky130_fd_pr__res_high_po_0p69 l=12.22
X28 a_6834_1206# a_6834_n1638# a_n7570_n1768# sky130_fd_pr__res_high_po_0p69 l=12.22
X29 a_n7440_1206# a_n7440_n1638# a_n7570_n1768# sky130_fd_pr__res_high_po_0p69 l=12.22
X30 a_750_1206# a_750_n1638# a_n7570_n1768# sky130_fd_pr__res_high_po_0p69 l=12.22
X31 a_2856_1206# a_2856_n1638# a_n7570_n1768# sky130_fd_pr__res_high_po_0p69 l=12.22
X32 a_n1122_1206# a_n1122_n1638# a_n7570_n1768# sky130_fd_pr__res_high_po_0p69 l=12.22
X33 a_4260_1206# a_4260_n1638# a_n7570_n1768# sky130_fd_pr__res_high_po_0p69 l=12.22
X34 a_n888_1206# a_n888_n1638# a_n7570_n1768# sky130_fd_pr__res_high_po_0p69 l=12.22
X35 a_n7206_1206# a_n7206_n1638# a_n7570_n1768# sky130_fd_pr__res_high_po_0p69 l=12.22
X36 a_n3228_1206# a_n3228_n1638# a_n7570_n1768# sky130_fd_pr__res_high_po_0p69 l=12.22
X37 a_2622_1206# a_2622_n1638# a_n7570_n1768# sky130_fd_pr__res_high_po_0p69 l=12.22
X38 a_6366_1206# a_6366_n1638# a_n7570_n1768# sky130_fd_pr__res_high_po_0p69 l=12.22
X39 a_6600_1206# a_6600_n1638# a_n7570_n1768# sky130_fd_pr__res_high_po_0p69 l=12.22
X40 a_282_1206# a_282_n1638# a_n7570_n1768# sky130_fd_pr__res_high_po_0p69 l=12.22
X41 a_2388_1206# a_2388_n1638# a_n7570_n1768# sky130_fd_pr__res_high_po_0p69 l=12.22
X42 a_n4866_1206# a_n4866_n1638# a_n7570_n1768# sky130_fd_pr__res_high_po_0p69 l=12.22
X43 a_4728_1206# a_4728_n1638# a_n7570_n1768# sky130_fd_pr__res_high_po_0p69 l=12.22
X44 a_n654_1206# a_n654_n1638# a_n7570_n1768# sky130_fd_pr__res_high_po_0p69 l=12.22
X45 a_n2292_1206# a_n2292_n1638# a_n7570_n1768# sky130_fd_pr__res_high_po_0p69 l=12.22
X46 a_2154_1206# a_2154_n1638# a_n7570_n1768# sky130_fd_pr__res_high_po_0p69 l=12.22
X47 a_6132_1206# a_6132_n1638# a_n7570_n1768# sky130_fd_pr__res_high_po_0p69 l=12.22
X48 a_n4632_1206# a_n4632_n1638# a_n7570_n1768# sky130_fd_pr__res_high_po_0p69 l=12.22
X49 a_n4398_1206# a_n4398_n1638# a_n7570_n1768# sky130_fd_pr__res_high_po_0p69 l=12.22
X50 a_3792_1206# a_3792_n1638# a_n7570_n1768# sky130_fd_pr__res_high_po_0p69 l=12.22
X51 a_n186_1206# a_n186_n1638# a_n7570_n1768# sky130_fd_pr__res_high_po_0p69 l=12.22
X52 a_n6738_1206# a_n6738_n1638# a_n7570_n1768# sky130_fd_pr__res_high_po_0p69 l=12.22
X53 a_n2760_1206# a_n2760_n1638# a_n7570_n1768# sky130_fd_pr__res_high_po_0p69 l=12.22
X54 a_516_1206# a_516_n1638# a_n7570_n1768# sky130_fd_pr__res_high_po_0p69 l=12.22
X55 a_5898_1206# a_5898_n1638# a_n7570_n1768# sky130_fd_pr__res_high_po_0p69 l=12.22
X56 a_n4164_1206# a_n4164_n1638# a_n7570_n1768# sky130_fd_pr__res_high_po_0p69 l=12.22
X57 a_4026_1206# a_4026_n1638# a_n7570_n1768# sky130_fd_pr__res_high_po_0p69 l=12.22
X58 a_n6504_1206# a_n6504_n1638# a_n7570_n1768# sky130_fd_pr__res_high_po_0p69 l=12.22
X59 a_n2526_1206# a_n2526_n1638# a_n7570_n1768# sky130_fd_pr__res_high_po_0p69 l=12.22
X60 a_1920_1206# a_1920_n1638# a_n7570_n1768# sky130_fd_pr__res_high_po_0p69 l=12.22
X61 a_n6270_1206# a_n6270_n1638# a_n7570_n1768# sky130_fd_pr__res_high_po_0p69 l=12.22
X62 a_1686_1206# a_1686_n1638# a_n7570_n1768# sky130_fd_pr__res_high_po_0p69 l=12.22
X63 a_5664_1206# a_5664_n1638# a_n7570_n1768# sky130_fd_pr__res_high_po_0p69 l=12.22
.ends

.subckt sky130_hcmus_ip__instramp VDD VSS G V1 V2 D0 D1 D2 D3 D4 D5 D6 D7 D8 D9 AVOUT1
+ AVOUT2 VOUT
Xx1 VDD x4/V2 D0 D3 D4 AVOUT1 D1 D2 G RB_array_20
Xx3 VDD x6/V2 D5 D8 D9 VOUT D6 D7 G RB_array_20
Xx2 VDD x5/V2 D0 D3 D4 AVOUT2 D1 D2 G RB_array_20
Xx4 V2 x4/V2 AVOUT1 VDD VSS opamp
Xx5 V1 x5/V2 AVOUT2 VDD VSS opamp
Xx6 x7/R1 x6/V2 VOUT VDD VSS opamp
XXR1 x4/V2 x5/V2 x5/V2 x4/V2 x4/V2 x5/V2 x4/V2 x5/V2 x5/V2 x5/V2 x4/V2 x5/V2 x4/V2
+ x5/V2 x4/V2 x4/V2 x5/V2 x5/V2 x5/V2 x4/V2 x4/V2 x5/V2 x5/V2 x4/V2 x5/V2 x5/V2 x5/V2
+ x4/V2 x4/V2 x4/V2 x4/V2 x4/V2 x5/V2 x5/V2 x4/V2 x5/V2 x5/V2 x5/V2 x4/V2 x5/V2 x4/V2
+ x5/V2 x4/V2 x5/V2 x4/V2 x4/V2 x5/V2 x5/V2 x4/V2 x5/V2 x4/V2 x4/V2 x4/V2 x4/V2 x5/V2
+ x4/V2 x5/V2 x5/V2 x4/V2 x5/V2 x5/V2 x5/V2 x4/V2 x4/V2 x5/V2 x5/V2 x4/V2 x5/V2 x4/V2
+ x4/V2 x4/V2 x5/V2 x5/V2 x4/V2 x5/V2 x5/V2 x5/V2 x4/V2 x4/V2 x4/V2 x4/V2 x5/V2 x5/V2
+ x4/V2 x4/V2 x4/V2 x5/V2 x4/V2 x5/V2 x4/V2 x5/V2 x4/V2 x4/V2 x4/V2 x4/V2 x5/V2 x5/V2
+ x4/V2 x4/V2 x4/V2 x5/V2 x5/V2 x4/V2 x5/V2 G x5/V2 x5/V2 x5/V2 x4/V2 x5/V2 x4/V2
+ x4/V2 x5/V2 x5/V2 x4/V2 x4/V2 x4/V2 x5/V2 x5/V2 x4/V2 x5/V2 x5/V2 x4/V2 x4/V2 x5/V2
+ x5/V2 x4/V2 x4/V2 x5/V2 sky130_fd_pr__res_high_po_0p69_WX3C5M
Xx7 VDD x7/R1 D5 D8 D9 G D6 D7 G RB_array_20
XXR2 x9/V2 x7/R1 x7/R1 x9/V2 x9/V2 x7/R1 x9/V2 x7/R1 x7/R1 x7/R1 x9/V2 x7/R1 x9/V2
+ x7/R1 x9/V2 x9/V2 x7/R1 x7/R1 x7/R1 x9/V2 x9/V2 x7/R1 x7/R1 x9/V2 x7/R1 x7/R1 x7/R1
+ x9/V2 x9/V2 x9/V2 x9/V2 x9/V2 x7/R1 x7/R1 x9/V2 x7/R1 x7/R1 x7/R1 x9/V2 x7/R1 x9/V2
+ x7/R1 x9/V2 x7/R1 x9/V2 x9/V2 x7/R1 x7/R1 x9/V2 x7/R1 x9/V2 x9/V2 x9/V2 x9/V2 x7/R1
+ x9/V2 x7/R1 x7/R1 x9/V2 x7/R1 x7/R1 x7/R1 x9/V2 x9/V2 x7/R1 x7/R1 x9/V2 x7/R1 x9/V2
+ x9/V2 x9/V2 x7/R1 x7/R1 x9/V2 x7/R1 x7/R1 x7/R1 x9/V2 x9/V2 x9/V2 x9/V2 x7/R1 x7/R1
+ x9/V2 x9/V2 x9/V2 x7/R1 x9/V2 x7/R1 x9/V2 x7/R1 x9/V2 x9/V2 x9/V2 x9/V2 x7/R1 x7/R1
+ x9/V2 x9/V2 x9/V2 x7/R1 x7/R1 x9/V2 x7/R1 G x7/R1 x7/R1 x7/R1 x9/V2 x7/R1 x9/V2
+ x9/V2 x7/R1 x7/R1 x9/V2 x9/V2 x9/V2 x7/R1 x7/R1 x9/V2 x7/R1 x7/R1 x9/V2 x9/V2 x7/R1
+ x7/R1 x9/V2 x9/V2 x7/R1 sky130_fd_pr__res_high_po_0p69_WX3C5M
Xx8 AVOUT1 x8/V2 x8/V2 VDD VSS opamp
Xx9 AVOUT2 x9/V2 x9/V2 VDD VSS opamp
XXR4 x8/V2 x6/V2 x6/V2 x8/V2 x8/V2 x6/V2 x8/V2 x6/V2 x6/V2 x6/V2 x8/V2 x6/V2 x8/V2
+ x6/V2 x8/V2 x8/V2 x6/V2 x6/V2 x6/V2 x8/V2 x8/V2 x6/V2 x6/V2 x8/V2 x6/V2 x6/V2 x6/V2
+ x8/V2 x8/V2 x8/V2 x8/V2 x8/V2 x6/V2 x6/V2 x8/V2 x6/V2 x6/V2 x6/V2 x8/V2 x6/V2 x8/V2
+ x6/V2 x8/V2 x6/V2 x8/V2 x8/V2 x6/V2 x6/V2 x8/V2 x6/V2 x8/V2 x8/V2 x8/V2 x8/V2 x6/V2
+ x8/V2 x6/V2 x6/V2 x8/V2 x6/V2 x6/V2 x6/V2 x8/V2 x8/V2 x6/V2 x6/V2 x8/V2 x6/V2 x8/V2
+ x8/V2 x8/V2 x6/V2 x6/V2 x8/V2 x6/V2 x6/V2 x6/V2 x8/V2 x8/V2 x8/V2 x8/V2 x6/V2 x6/V2
+ x8/V2 x8/V2 x8/V2 x6/V2 x8/V2 x6/V2 x8/V2 x6/V2 x8/V2 x8/V2 x8/V2 x8/V2 x6/V2 x6/V2
+ x8/V2 x8/V2 x8/V2 x6/V2 x6/V2 x8/V2 x6/V2 G x6/V2 x6/V2 x6/V2 x8/V2 x6/V2 x8/V2
+ x8/V2 x6/V2 x6/V2 x8/V2 x8/V2 x8/V2 x6/V2 x6/V2 x8/V2 x6/V2 x6/V2 x8/V2 x8/V2 x6/V2
+ x6/V2 x8/V2 x8/V2 x6/V2 sky130_fd_pr__res_high_po_0p69_WX3C5M
.ends

