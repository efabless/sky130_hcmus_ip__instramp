magic
tech sky130A
magscale 1 2
timestamp 1716807968
<< pwell >>
rect -328 -1167 328 1167
<< mvnmos >>
rect -100 109 100 909
rect -100 -909 100 -109
<< mvndiff >>
rect -158 897 -100 909
rect -158 121 -146 897
rect -112 121 -100 897
rect -158 109 -100 121
rect 100 897 158 909
rect 100 121 112 897
rect 146 121 158 897
rect 100 109 158 121
rect -158 -121 -100 -109
rect -158 -897 -146 -121
rect -112 -897 -100 -121
rect -158 -909 -100 -897
rect 100 -121 158 -109
rect 100 -897 112 -121
rect 146 -897 158 -121
rect 100 -909 158 -897
<< mvndiffc >>
rect -146 121 -112 897
rect 112 121 146 897
rect -146 -897 -112 -121
rect 112 -897 146 -121
<< mvpsubdiff >>
rect -292 1119 292 1131
rect -292 1085 -184 1119
rect 184 1085 292 1119
rect -292 1073 292 1085
rect -292 1023 -234 1073
rect -292 -1023 -280 1023
rect -246 -1023 -234 1023
rect 234 1023 292 1073
rect -292 -1073 -234 -1023
rect 234 -1023 246 1023
rect 280 -1023 292 1023
rect 234 -1073 292 -1023
rect -292 -1085 292 -1073
rect -292 -1119 -184 -1085
rect 184 -1119 292 -1085
rect -292 -1131 292 -1119
<< mvpsubdiffcont >>
rect -184 1085 184 1119
rect -280 -1023 -246 1023
rect 246 -1023 280 1023
rect -184 -1119 184 -1085
<< poly >>
rect -100 981 100 997
rect -100 947 -84 981
rect 84 947 100 981
rect -100 909 100 947
rect -100 71 100 109
rect -100 37 -84 71
rect 84 37 100 71
rect -100 21 100 37
rect -100 -37 100 -21
rect -100 -71 -84 -37
rect 84 -71 100 -37
rect -100 -109 100 -71
rect -100 -947 100 -909
rect -100 -981 -84 -947
rect 84 -981 100 -947
rect -100 -997 100 -981
<< polycont >>
rect -84 947 84 981
rect -84 37 84 71
rect -84 -71 84 -37
rect -84 -981 84 -947
<< locali >>
rect -280 1085 -184 1119
rect 184 1085 280 1119
rect -280 1023 -246 1085
rect 246 1023 280 1085
rect -100 947 -84 981
rect 84 947 100 981
rect -146 897 -112 913
rect -146 105 -112 121
rect 112 897 146 913
rect 112 105 146 121
rect -100 37 -84 71
rect 84 37 100 71
rect -100 -71 -84 -37
rect 84 -71 100 -37
rect -146 -121 -112 -105
rect -146 -913 -112 -897
rect 112 -121 146 -105
rect 112 -913 146 -897
rect -100 -981 -84 -947
rect 84 -981 100 -947
rect -280 -1085 -246 -1023
rect 246 -1085 280 -1023
rect -280 -1119 -184 -1085
rect 184 -1119 280 -1085
<< viali >>
rect -84 947 84 981
rect -146 121 -112 897
rect 112 121 146 897
rect -84 37 84 71
rect -84 -71 84 -37
rect -146 -897 -112 -121
rect 112 -897 146 -121
rect -84 -981 84 -947
<< metal1 >>
rect -96 981 96 987
rect -96 947 -84 981
rect 84 947 96 981
rect -96 941 96 947
rect -152 897 -106 909
rect -152 121 -146 897
rect -112 121 -106 897
rect -152 109 -106 121
rect 106 897 152 909
rect 106 121 112 897
rect 146 121 152 897
rect 106 109 152 121
rect -96 71 96 77
rect -96 37 -84 71
rect 84 37 96 71
rect -96 31 96 37
rect -96 -37 96 -31
rect -96 -71 -84 -37
rect 84 -71 96 -37
rect -96 -77 96 -71
rect -152 -121 -106 -109
rect -152 -897 -146 -121
rect -112 -897 -106 -121
rect -152 -909 -106 -897
rect 106 -121 152 -109
rect 106 -897 112 -121
rect 146 -897 152 -121
rect 106 -909 152 -897
rect -96 -947 96 -941
rect -96 -981 -84 -947
rect 84 -981 96 -947
rect -96 -987 96 -981
<< properties >>
string FIXED_BBOX -263 -1102 263 1102
string gencell sky130_fd_pr__nfet_g5v0d10v5
string library sky130
string parameters w 4.0 l 1.0 m 2 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
