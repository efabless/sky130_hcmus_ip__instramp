magic
tech sky130A
magscale 1 2
timestamp 1716789169
<< nwell >>
rect -745 -2126 745 2126
<< mvpmos >>
rect -487 -1900 -287 1900
rect -229 -1900 -29 1900
rect 29 -1900 229 1900
rect 287 -1900 487 1900
<< mvpdiff >>
rect -545 1888 -487 1900
rect -545 -1888 -533 1888
rect -499 -1888 -487 1888
rect -545 -1900 -487 -1888
rect -287 1888 -229 1900
rect -287 -1888 -275 1888
rect -241 -1888 -229 1888
rect -287 -1900 -229 -1888
rect -29 1888 29 1900
rect -29 -1888 -17 1888
rect 17 -1888 29 1888
rect -29 -1900 29 -1888
rect 229 1888 287 1900
rect 229 -1888 241 1888
rect 275 -1888 287 1888
rect 229 -1900 287 -1888
rect 487 1888 545 1900
rect 487 -1888 499 1888
rect 533 -1888 545 1888
rect 487 -1900 545 -1888
<< mvpdiffc >>
rect -533 -1888 -499 1888
rect -275 -1888 -241 1888
rect -17 -1888 17 1888
rect 241 -1888 275 1888
rect 499 -1888 533 1888
<< mvnsubdiff >>
rect -679 2048 679 2060
rect -679 2014 -571 2048
rect 571 2014 679 2048
rect -679 2002 679 2014
rect -679 1952 -621 2002
rect -679 -1952 -667 1952
rect -633 -1952 -621 1952
rect 621 1952 679 2002
rect -679 -2002 -621 -1952
rect 621 -1952 633 1952
rect 667 -1952 679 1952
rect 621 -2002 679 -1952
rect -679 -2014 679 -2002
rect -679 -2048 -571 -2014
rect 571 -2048 679 -2014
rect -679 -2060 679 -2048
<< mvnsubdiffcont >>
rect -571 2014 571 2048
rect -667 -1952 -633 1952
rect 633 -1952 667 1952
rect -571 -2048 571 -2014
<< poly >>
rect -487 1900 -287 1926
rect -229 1900 -29 1926
rect 29 1900 229 1926
rect 287 1900 487 1926
rect -487 -1926 -287 -1900
rect -229 -1926 -29 -1900
rect 29 -1926 229 -1900
rect 287 -1926 487 -1900
<< locali >>
rect -667 2014 -571 2048
rect 571 2014 667 2048
rect -667 1952 -633 2014
rect 633 1952 667 2014
rect -533 1888 -499 1904
rect -533 -1904 -499 -1888
rect -275 1888 -241 1904
rect -275 -1904 -241 -1888
rect -17 1888 17 1904
rect -17 -1904 17 -1888
rect 241 1888 275 1904
rect 241 -1904 275 -1888
rect 499 1888 533 1904
rect 499 -1904 533 -1888
rect -667 -2014 -633 -1952
rect 633 -2014 667 -1952
rect -667 -2048 -571 -2014
rect 571 -2048 667 -2014
<< viali >>
rect -533 -1888 -499 1888
rect -275 -1888 -241 1888
rect -17 -1888 17 1888
rect 241 -1888 275 1888
rect 499 -1888 533 1888
<< metal1 >>
rect -539 1888 -493 1900
rect -539 -1888 -533 1888
rect -499 -1888 -493 1888
rect -539 -1900 -493 -1888
rect -281 1888 -235 1900
rect -281 -1888 -275 1888
rect -241 -1888 -235 1888
rect -281 -1900 -235 -1888
rect -23 1888 23 1900
rect -23 -1888 -17 1888
rect 17 -1888 23 1888
rect -23 -1900 23 -1888
rect 235 1888 281 1900
rect 235 -1888 241 1888
rect 275 -1888 281 1888
rect 235 -1900 281 -1888
rect 493 1888 539 1900
rect 493 -1888 499 1888
rect 533 -1888 539 1888
rect 493 -1900 539 -1888
<< properties >>
string FIXED_BBOX -650 -2031 650 2031
string gencell sky130_fd_pr__pfet_g5v0d10v5
string library sky130
string parameters w 19.0 l 1.0 m 1 nf 4 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 0 botc 0 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
