magic
tech sky130A
magscale 1 2
timestamp 1720369107
<< locali >>
rect 2065 16111 3639 16253
rect 2065 15773 2207 16111
rect 3497 15776 3639 16111
rect 2065 15760 2220 15773
rect 2065 14973 2144 15760
rect 2186 14973 2220 15760
rect 2065 14949 2220 14973
rect 3482 15757 3639 15776
rect 3482 14970 3511 15757
rect 3553 14970 3639 15757
rect 3482 14952 3639 14970
rect -53 13228 1057 13392
rect -53 12635 111 13228
rect 893 12635 1057 13228
rect 2065 12645 2207 14949
rect 3497 12654 3639 14952
rect -53 12599 1057 12635
rect -53 12574 1061 12599
rect -53 12441 3623 12574
rect -53 12090 111 12441
rect 893 12435 3623 12441
rect -53 11330 -36 12090
rect 95 11330 111 12090
rect -53 8998 111 11330
rect 3459 12089 3623 12435
rect 3459 11329 3472 12089
rect 3603 11329 3623 12089
rect 3459 9000 3623 11329
<< viali >>
rect 2144 14973 2186 15760
rect 3511 14970 3553 15757
rect -36 11330 95 12090
rect 3472 11329 3603 12089
<< metal1 >>
rect 2401 16331 3287 16335
rect 2401 16260 2421 16331
rect 2717 16260 3287 16331
rect 2401 16254 3287 16260
rect 2415 15983 2496 16254
rect 3206 15987 3287 16254
rect 2415 15979 2501 15983
rect 2117 15763 2220 15773
rect 2117 14970 2131 15763
rect 2210 14970 2220 15763
rect 2117 14949 2220 14970
rect 2288 14827 2381 14855
rect 177 13010 283 13020
rect 177 12835 197 13010
rect 260 12835 283 13010
rect 177 12781 283 12835
rect 328 12781 404 13099
rect 441 13010 547 13023
rect 441 12835 464 13010
rect 527 12835 547 13010
rect 441 12824 547 12835
rect 441 12781 547 12782
rect 586 12781 662 13099
rect 698 13010 804 13027
rect 698 12835 718 13010
rect 781 12835 804 13010
rect 2288 12911 2301 14827
rect 2369 12911 2381 14827
rect 2288 12882 2381 12911
rect 698 12781 804 12835
rect 2433 12784 2501 15979
rect 2554 12841 2629 14841
rect 177 12736 804 12781
rect 267 12735 717 12736
rect 328 12572 404 12735
rect 586 12572 662 12735
rect 2679 12709 2747 15972
rect 2807 15895 2900 15911
rect 2807 12890 2828 15895
rect 2884 12890 2900 15895
rect 2807 12864 2900 12890
rect 2953 12913 3021 15979
rect 3070 12913 3145 14830
rect 2953 12843 3145 12913
rect 2953 12791 3021 12843
rect 3070 12841 3145 12843
rect 2952 12780 3021 12791
rect 2952 12709 3020 12780
rect 3202 12777 3270 15976
rect 3482 15757 3585 15776
rect 3482 15755 3511 15757
rect 3553 15755 3585 15757
rect 3482 14962 3490 15755
rect 3569 14962 3585 15755
rect 3482 14952 3585 14962
rect 3319 14825 3412 14853
rect 3319 12909 3332 14825
rect 3400 12909 3412 14825
rect 3319 12880 3412 12909
rect 2679 12641 3020 12709
rect 328 12535 3240 12572
rect 328 12473 3242 12535
rect -53 12090 116 12108
rect 210 12092 216 12138
rect 250 12092 256 12138
rect -53 11330 -36 12090
rect 95 11330 116 12090
rect -53 11311 116 11330
rect 191 12084 273 12092
rect 191 10324 197 12084
rect 268 10324 273 12084
rect 191 9347 273 10324
rect 210 9332 216 9347
rect 250 9332 256 9347
rect 328 9154 404 12473
rect 449 11152 531 12092
rect 449 9380 455 11152
rect 526 9380 531 11152
rect 449 9347 531 9380
rect 586 9154 662 12473
rect 726 12092 732 12120
rect 766 12092 772 12120
rect 707 12084 789 12092
rect 707 10324 713 12084
rect 784 10324 789 12084
rect 707 9361 789 10324
rect 844 9154 920 12473
rect 984 12092 990 12120
rect 1024 12092 1030 12120
rect 965 11152 1047 12092
rect 965 9380 971 11152
rect 1042 9380 1047 11152
rect 965 9361 1047 9380
rect 1102 9154 1178 12473
rect 1242 12092 1248 12120
rect 1282 12092 1288 12120
rect 1223 12084 1305 12092
rect 1223 10324 1229 12084
rect 1300 10324 1305 12084
rect 1223 9361 1305 10324
rect 1360 9154 1436 12473
rect 1500 12092 1506 12120
rect 1540 12092 1546 12120
rect 1481 11152 1563 12092
rect 1481 9380 1487 11152
rect 1558 9380 1563 11152
rect 1481 9361 1563 9380
rect 1618 9154 1694 12473
rect 1758 12092 1764 12120
rect 1798 12092 1804 12120
rect 1739 12084 1821 12092
rect 1739 10324 1745 12084
rect 1816 10324 1821 12084
rect 1739 9361 1821 10324
rect 1876 9154 1952 12473
rect 2016 12092 2022 12120
rect 2056 12092 2062 12120
rect 1997 11152 2079 12092
rect 1997 9380 2003 11152
rect 2074 9380 2079 11152
rect 1997 9361 2079 9380
rect 2134 9154 2210 12473
rect 2274 12092 2280 12120
rect 2314 12092 2320 12120
rect 2255 12084 2337 12092
rect 2255 10324 2261 12084
rect 2332 10324 2337 12084
rect 2255 9361 2337 10324
rect 2392 9154 2468 12473
rect 2532 12092 2538 12120
rect 2572 12092 2578 12120
rect 2513 11152 2595 12092
rect 2513 9380 2519 11152
rect 2590 9380 2595 11152
rect 2513 9361 2595 9380
rect 2650 9154 2726 12473
rect 2790 12092 2796 12120
rect 2830 12092 2836 12120
rect 2771 12084 2853 12092
rect 2771 10324 2777 12084
rect 2848 10324 2853 12084
rect 2771 9361 2853 10324
rect 2908 9154 2984 12473
rect 3048 12092 3054 12120
rect 3088 12092 3094 12120
rect 3029 11152 3111 12092
rect 3029 9380 3035 11152
rect 3106 9380 3111 11152
rect 3029 9361 3111 9380
rect 3166 9154 3242 12473
rect 3306 12092 3312 12120
rect 3346 12092 3352 12120
rect 3287 12084 3369 12092
rect 3287 10324 3293 12084
rect 3364 10324 3369 12084
rect 3455 12089 3624 12107
rect 3455 11329 3472 12089
rect 3603 11329 3624 12089
rect 3455 11310 3624 11329
rect 3287 9361 3369 10324
<< via1 >>
rect 2421 16260 2717 16331
rect 2131 15760 2210 15763
rect 2131 14973 2144 15760
rect 2144 14973 2186 15760
rect 2186 14973 2210 15760
rect 2131 14970 2210 14973
rect 197 12835 260 13010
rect 464 12835 527 13010
rect 718 12835 781 13010
rect 2301 12911 2369 14827
rect 2828 12890 2884 15895
rect 3490 14970 3511 15755
rect 3511 14970 3553 15755
rect 3553 14970 3569 15755
rect 3490 14962 3569 14970
rect 3332 12909 3400 14825
rect -36 11330 95 12090
rect 197 10324 268 12084
rect 455 9380 526 11152
rect 713 10324 784 12084
rect 971 9380 1042 11152
rect 1229 10324 1300 12084
rect 1487 9380 1558 11152
rect 1745 10324 1816 12084
rect 2003 9380 2074 11152
rect 2261 10324 2332 12084
rect 2519 9380 2590 11152
rect 2777 10324 2848 12084
rect 3035 9380 3106 11152
rect 3293 10324 3364 12084
rect 3472 11329 3603 12089
<< metal2 >>
rect 2401 16331 2736 16335
rect 2401 16322 2421 16331
rect -108 16266 2421 16322
rect 2401 16260 2421 16266
rect 2717 16260 2736 16331
rect 2401 16254 2736 16260
rect 2807 15895 2900 15911
rect 2807 15783 2828 15895
rect -108 15763 2828 15783
rect -108 14970 2131 15763
rect 2210 14970 2828 15763
rect -108 14936 2828 14970
rect 2253 14827 2404 14859
rect 2253 13293 2301 14827
rect 177 13126 2301 13293
rect 177 13010 283 13126
rect 177 12835 197 13010
rect 260 12835 283 13010
rect 177 12819 283 12835
rect 393 13010 599 13023
rect 393 12835 464 13010
rect 527 12835 599 13010
rect 393 12107 599 12835
rect 698 13010 804 13126
rect 698 12835 718 13010
rect 781 12835 804 13010
rect 2253 12911 2301 13126
rect 2369 12911 2404 14827
rect 2253 12886 2404 12911
rect 2565 12890 2828 14936
rect 2884 15783 2900 15895
rect 2884 15755 3589 15783
rect 2884 14962 3490 15755
rect 3569 14962 3589 15755
rect 2884 14936 3589 14962
rect 2884 12890 3141 14936
rect 3319 14849 3412 14853
rect 2288 12882 2381 12886
rect 2565 12865 3141 12890
rect 3296 14847 3447 14849
rect 3754 14847 3945 16552
rect 3296 14825 3945 14847
rect 3296 12909 3332 14825
rect 3400 14656 3945 14825
rect 3400 12909 3447 14656
rect 3296 12876 3447 12909
rect 2807 12864 2900 12865
rect 698 12826 804 12835
rect -108 12090 3657 12107
rect -108 11330 -36 12090
rect 95 12089 3657 12090
rect 95 12084 3472 12089
rect 95 11330 197 12084
rect -108 11310 197 11330
rect 268 11310 713 12084
rect 197 10311 268 10324
rect 419 11152 541 11183
rect 419 9380 455 11152
rect 526 9380 541 11152
rect 784 11310 1229 12084
rect 713 10311 784 10324
rect 935 11152 1057 11183
rect 419 9302 541 9380
rect 935 9380 971 11152
rect 1042 9380 1057 11152
rect 1300 11310 1745 12084
rect 1229 10311 1300 10324
rect 1451 11152 1573 11183
rect 935 9302 1057 9380
rect 1451 9380 1487 11152
rect 1558 9380 1573 11152
rect 1816 11310 2261 12084
rect 1745 10311 1816 10324
rect 1967 11152 2089 11183
rect 1451 9302 1573 9380
rect 1967 9380 2003 11152
rect 2074 9380 2089 11152
rect 2332 11310 2777 12084
rect 2261 10311 2332 10324
rect 2483 11152 2605 11183
rect 1967 9302 2089 9380
rect 2483 9847 2519 11152
rect 2590 9847 2605 11152
rect 2848 11310 3293 12084
rect 2777 10311 2848 10324
rect 2999 11152 3121 11183
rect 2483 9321 2494 9847
rect 2594 9321 2605 9847
rect 2483 9302 2605 9321
rect 2999 10039 3035 11152
rect 3106 10039 3121 11152
rect 3364 11329 3472 12084
rect 3603 11329 3657 12089
rect 3364 11310 3657 11329
rect 3293 10311 3364 10324
rect 2999 9465 3009 10039
rect 3109 9465 3121 10039
rect 2999 9380 3035 9465
rect 3106 9380 3121 9465
rect 2999 9302 3121 9380
rect 444 8952 515 9302
rect 957 8952 1028 9302
rect 1475 9061 1546 9302
rect 1995 9226 2066 9302
rect 1995 9155 4002 9226
rect 1475 8990 4002 9061
<< via2 >>
rect 2494 9380 2519 9847
rect 2519 9380 2590 9847
rect 2590 9380 2594 9847
rect 2494 9321 2594 9380
rect 3009 9465 3035 10039
rect 3035 9465 3106 10039
rect 3106 9465 3109 10039
<< metal3 >>
rect 3000 10039 3120 10051
rect 2485 9847 2605 9862
rect 2485 9321 2494 9847
rect 2594 9341 2605 9847
rect 3000 9465 3009 10039
rect 3109 9531 3120 10039
rect 3109 9465 4002 9531
rect 3000 9452 4002 9465
rect 3000 9451 3120 9452
rect 2594 9321 4002 9341
rect 2485 9262 4002 9321
use sky130_fd_pr__nfet_g5v0d10v5_EHZ5KL  sky130_fd_pr__nfet_g5v0d10v5_EHZ5KL_0 paramcells
timestamp 1720214482
transform 1 0 2851 0 1 14380
box -715 -1802 715 1802
use sky130_fd_pr__pfet_g5v0d10v5_6HDYS4  sky130_fd_pr__pfet_g5v0d10v5_6HDYS4_0 paramcells
timestamp 1720214482
transform 1 0 491 0 1 12923
box -487 -397 487 397
use sky130_fd_pr__pfet_g5v0d10v5_SKQKSC  sky130_fd_pr__pfet_g5v0d10v5_SKQKSC_0 paramcells
timestamp 1720214482
transform -1 0 1781 0 -1 10729
box -1777 -1797 1777 1797
<< labels >>
flabel metal2 3754 16382 3945 16552 0 FreeSans 960 90 0 0 ibias
port 0 nsew
flabel metal2 -108 14936 141 15783 0 FreeSans 1600 90 0 0 VSS
port 1 nsew
flabel metal2 -108 11310 -36 12107 0 FreeSans 1600 90 0 0 VDD
port 2 nsew
flabel metal2 -108 16266 58 16322 0 FreeSans 960 0 0 0 ena3v3
port 3 nsew
flabel metal2 444 8952 515 9101 0 FreeSans 960 90 0 0 ibias0
port 4 nsew
flabel metal2 957 8952 1028 9101 0 FreeSans 960 90 0 0 ibias1
port 5 nsew
flabel metal2 3849 8990 4002 9061 0 FreeSans 960 0 0 0 ibias2
port 6 nsew
flabel metal2 3849 9155 4002 9226 0 FreeSans 960 0 0 0 ibias3
port 7 nsew
flabel metal3 3842 9262 4002 9341 0 FreeSans 960 0 0 0 ibias4
port 8 nsew
flabel metal3 3842 9452 4002 9531 0 FreeSans 960 0 0 0 ibias5
port 9 nsew
<< end >>
