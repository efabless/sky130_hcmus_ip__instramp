magic
tech sky130A
magscale 1 2
timestamp 1720214482
<< pwell >>
rect -715 -1802 715 1802
<< mvnmos >>
rect -487 -1544 -287 1544
rect -229 -1544 -29 1544
rect 29 -1544 229 1544
rect 287 -1544 487 1544
<< mvndiff >>
rect -545 1532 -487 1544
rect -545 -1532 -533 1532
rect -499 -1532 -487 1532
rect -545 -1544 -487 -1532
rect -287 1532 -229 1544
rect -287 -1532 -275 1532
rect -241 -1532 -229 1532
rect -287 -1544 -229 -1532
rect -29 1532 29 1544
rect -29 -1532 -17 1532
rect 17 -1532 29 1532
rect -29 -1544 29 -1532
rect 229 1532 287 1544
rect 229 -1532 241 1532
rect 275 -1532 287 1532
rect 229 -1544 287 -1532
rect 487 1532 545 1544
rect 487 -1532 499 1532
rect 533 -1532 545 1532
rect 487 -1544 545 -1532
<< mvndiffc >>
rect -533 -1532 -499 1532
rect -275 -1532 -241 1532
rect -17 -1532 17 1532
rect 241 -1532 275 1532
rect 499 -1532 533 1532
<< mvpsubdiff >>
rect -679 1754 679 1766
rect -679 1720 -571 1754
rect 571 1720 679 1754
rect -679 1708 679 1720
rect -679 1658 -621 1708
rect -679 -1658 -667 1658
rect -633 -1658 -621 1658
rect 621 1658 679 1708
rect -679 -1708 -621 -1658
rect 621 -1658 633 1658
rect 667 -1658 679 1658
rect 621 -1708 679 -1658
rect -679 -1720 679 -1708
rect -679 -1754 -571 -1720
rect 571 -1754 679 -1720
rect -679 -1766 679 -1754
<< mvpsubdiffcont >>
rect -571 1720 571 1754
rect -667 -1658 -633 1658
rect 633 -1658 667 1658
rect -571 -1754 571 -1720
<< poly >>
rect -487 1616 -287 1632
rect -487 1582 -471 1616
rect -303 1582 -287 1616
rect -487 1544 -287 1582
rect -229 1616 -29 1632
rect -229 1582 -213 1616
rect -45 1582 -29 1616
rect -229 1544 -29 1582
rect 29 1616 229 1632
rect 29 1582 45 1616
rect 213 1582 229 1616
rect 29 1544 229 1582
rect 287 1616 487 1632
rect 287 1582 303 1616
rect 471 1582 487 1616
rect 287 1544 487 1582
rect -487 -1582 -287 -1544
rect -487 -1616 -471 -1582
rect -303 -1616 -287 -1582
rect -487 -1632 -287 -1616
rect -229 -1582 -29 -1544
rect -229 -1616 -213 -1582
rect -45 -1616 -29 -1582
rect -229 -1632 -29 -1616
rect 29 -1582 229 -1544
rect 29 -1616 45 -1582
rect 213 -1616 229 -1582
rect 29 -1632 229 -1616
rect 287 -1582 487 -1544
rect 287 -1616 303 -1582
rect 471 -1616 487 -1582
rect 287 -1632 487 -1616
<< polycont >>
rect -471 1582 -303 1616
rect -213 1582 -45 1616
rect 45 1582 213 1616
rect 303 1582 471 1616
rect -471 -1616 -303 -1582
rect -213 -1616 -45 -1582
rect 45 -1616 213 -1582
rect 303 -1616 471 -1582
<< locali >>
rect -667 1720 -571 1754
rect 571 1720 667 1754
rect -667 1658 -633 1720
rect 633 1658 667 1720
rect -487 1582 -471 1616
rect -303 1582 -287 1616
rect -229 1582 -213 1616
rect -45 1582 -29 1616
rect 29 1582 45 1616
rect 213 1582 229 1616
rect 287 1582 303 1616
rect 471 1582 487 1616
rect -533 1532 -499 1548
rect -533 -1548 -499 -1532
rect -275 1532 -241 1548
rect -275 -1548 -241 -1532
rect -17 1532 17 1548
rect -17 -1548 17 -1532
rect 241 1532 275 1548
rect 241 -1548 275 -1532
rect 499 1532 533 1548
rect 499 -1548 533 -1532
rect -487 -1616 -471 -1582
rect -303 -1616 -287 -1582
rect -229 -1616 -213 -1582
rect -45 -1616 -29 -1582
rect 29 -1616 45 -1582
rect 213 -1616 229 -1582
rect 287 -1616 303 -1582
rect 471 -1616 487 -1582
rect -667 -1720 -633 -1658
rect 633 -1720 667 -1658
rect -667 -1754 -571 -1720
rect 571 -1754 667 -1720
<< viali >>
rect -471 1582 -303 1616
rect -213 1582 -45 1616
rect 45 1582 213 1616
rect 303 1582 471 1616
rect -533 -1532 -499 1532
rect -275 -1532 -241 1532
rect -17 -1532 17 1532
rect 241 -1532 275 1532
rect 499 -1532 533 1532
rect -471 -1616 -303 -1582
rect -213 -1616 -45 -1582
rect 45 -1616 213 -1582
rect 303 -1616 471 -1582
<< metal1 >>
rect -483 1616 -291 1622
rect -483 1582 -471 1616
rect -303 1582 -291 1616
rect -483 1576 -291 1582
rect -225 1616 -33 1622
rect -225 1582 -213 1616
rect -45 1582 -33 1616
rect -225 1576 -33 1582
rect 33 1616 225 1622
rect 33 1582 45 1616
rect 213 1582 225 1616
rect 33 1576 225 1582
rect 291 1616 483 1622
rect 291 1582 303 1616
rect 471 1582 483 1616
rect 291 1576 483 1582
rect -539 1532 -493 1544
rect -539 -1532 -533 1532
rect -499 -1532 -493 1532
rect -539 -1544 -493 -1532
rect -281 1532 -235 1544
rect -281 -1532 -275 1532
rect -241 -1532 -235 1532
rect -281 -1544 -235 -1532
rect -23 1532 23 1544
rect -23 -1532 -17 1532
rect 17 -1532 23 1532
rect -23 -1544 23 -1532
rect 235 1532 281 1544
rect 235 -1532 241 1532
rect 275 -1532 281 1532
rect 235 -1544 281 -1532
rect 493 1532 539 1544
rect 493 -1532 499 1532
rect 533 -1532 539 1532
rect 493 -1544 539 -1532
rect -483 -1582 -291 -1576
rect -483 -1616 -471 -1582
rect -303 -1616 -291 -1582
rect -483 -1622 -291 -1616
rect -225 -1582 -33 -1576
rect -225 -1616 -213 -1582
rect -45 -1616 -33 -1582
rect -225 -1622 -33 -1616
rect 33 -1582 225 -1576
rect 33 -1616 45 -1582
rect 213 -1616 225 -1582
rect 33 -1622 225 -1616
rect 291 -1582 483 -1576
rect 291 -1616 303 -1582
rect 471 -1616 483 -1582
rect 291 -1622 483 -1616
<< properties >>
string FIXED_BBOX -650 -1737 650 1737
string gencell sky130_fd_pr__nfet_g5v0d10v5
string library sky130
string parameters w 15.44 l 1 m 1 nf 4 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
