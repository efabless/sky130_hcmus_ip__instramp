magic
tech sky130A
magscale 1 2
timestamp 1716878682
<< error_s >>
rect 763 4032 798 4066
rect 764 4013 798 4032
rect 783 530 798 4013
rect 817 3979 852 4013
rect 1180 3979 1215 4013
rect 817 530 851 3979
rect 1181 3960 1215 3979
rect 817 496 832 530
rect 1200 477 1215 3960
rect 1234 3926 1269 3960
rect 1234 477 1268 3926
rect 1234 443 1249 477
rect 3010 253 3057 1497
rect 3064 199 3111 1551
rect 3601 188 3648 2450
rect 3655 134 3702 2504
use sky130_fd_pr__nfet_g5v0d10v5_KE4BRS  XM1
timestamp 1716807968
transform 1 0 6698 0 1 896
box -715 -1069 715 1069
use sky130_fd_pr__nfet_g5v0d10v5_WVAQGW  XM6
timestamp 1716807968
transform 1 0 2765 0 1 875
box -328 -658 328 658
use sky130_fd_pr__nfet_g5v0d10v5_MMMQGW  XM7
timestamp 1716807968
transform 1 0 3356 0 1 1319
box -328 -1167 328 1167
use sky130_fd_pr__nfet_g5v0d10v5_FVDQGW  XM8
timestamp 1716807968
transform 1 0 3947 0 1 2272
box -328 -2185 328 2185
use sky130_fd_pr__nfet_g5v0d10v5_KVPNGW  XM9
timestamp 1716807968
transform 1 0 6350 0 1 8023
box -328 -4221 328 4221
use sky130_fd_pr__nfet_g5v0d10v5_NEKL4L  XM10
timestamp 1716878682
transform 1 0 10640 0 1 13085
box -158 -8919 158 8919
use sky130_fd_pr__nfet_g5v0d10v5_DX5ZG7  XM11
timestamp 1716807968
transform 1 0 5318 0 1 1073
box -328 -1385 328 1385
use sky130_fd_pr__res_high_po_0p69_JKKHRG  XR1
timestamp 1716807968
transform 1 0 599 0 1 2298
box -235 -1804 235 1804
use sky130_fd_pr__res_high_po_0p69_JKKHRG  XR2
timestamp 1716807968
transform 1 0 -1663 0 1 2450
box -235 -1804 235 1804
use sky130_fd_pr__res_high_po_0p69_JKKHRG  XR3
timestamp 1716807968
transform 1 0 1016 0 1 2245
box -235 -1804 235 1804
use sky130_fd_pr__res_high_po_0p69_JKKHRG  XR4
timestamp 1716807968
transform 1 0 1433 0 1 2192
box -235 -1804 235 1804
use sky130_fd_pr__res_high_po_0p69_JKKHRG  XR5
timestamp 1716807968
transform 1 0 -6165 0 1 2052
box -235 -1804 235 1804
use sky130_fd_pr__res_high_po_0p69_HBQF5Z  XR6
timestamp 1716807968
transform 1 0 1658 0 1 6596
box -1990 -1804 1990 1804
<< end >>
