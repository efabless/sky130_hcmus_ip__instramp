* SPICE3 file created from opamp.ext - technology: sky130A

.subckt sky130_fd_pr__res_high_po_0p69_T8KQH6 a_n199_n866# a_n69_n736# a_n69_304#
X0 a_n69_304# a_n69_n736# a_n199_n866# sky130_fd_pr__res_high_po_0p69 l=3.04
C0 a_n69_304# a_n69_n736# 0.0134f
C1 a_n69_n736# a_n199_n866# 0.659f
C2 a_n69_304# a_n199_n866# 0.659f
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_K8DQNF a_n29_n1536# a_229_n1536# a_n229_n1562#
+ w_n487_n1762# a_n287_n1536# a_29_n1562# VSUBS
X0 a_n29_n1536# a_n229_n1562# a_n287_n1536# w_n487_n1762# sky130_fd_pr__pfet_g5v0d10v5 ad=2.17 pd=15.3 as=4.35 ps=30.6 w=15 l=1
X1 a_229_n1536# a_29_n1562# a_n29_n1536# w_n487_n1762# sky130_fd_pr__pfet_g5v0d10v5 ad=4.35 pd=30.6 as=2.17 ps=15.3 w=15 l=1
C0 a_229_n1536# a_29_n1562# 0.326f
C1 w_n487_n1762# a_n29_n1536# 0.023f
C2 w_n487_n1762# a_n287_n1536# 0.868f
C3 a_n29_n1536# a_n229_n1562# 0.326f
C4 a_n287_n1536# a_n229_n1562# 0.326f
C5 a_n29_n1536# a_29_n1562# 0.326f
C6 w_n487_n1762# a_n229_n1562# 0.257f
C7 a_n29_n1536# a_229_n1536# 0.82f
C8 w_n487_n1762# a_29_n1562# 0.257f
C9 a_29_n1562# a_n229_n1562# 0.0619f
C10 w_n487_n1762# a_229_n1536# 0.868f
C11 a_n287_n1536# a_n29_n1536# 0.82f
C12 a_229_n1536# VSUBS 0.733f
C13 a_n29_n1536# VSUBS 0.418f
C14 a_n287_n1536# VSUBS 0.733f
C15 a_29_n1562# VSUBS 0.228f
C16 a_n229_n1562# VSUBS 0.228f
C17 w_n487_n1762# VSUBS 12.4f
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_VYCZE8 a_100_n1681# a_n292_n1841# a_n100_n1707#
+ a_n158_n1681#
X0 a_100_n1681# a_n100_n1707# a_n158_n1681# a_n292_n1841# sky130_fd_pr__nfet_g5v0d10v5 ad=4.78 pd=33.6 as=4.78 ps=33.6 w=16.5 l=1
C0 a_n100_n1707# a_n158_n1681# 0.358f
C1 a_n100_n1707# a_100_n1681# 0.358f
C2 a_100_n1681# a_n158_n1681# 0.901f
C3 a_100_n1681# a_n292_n1841# 1.75f
C4 a_n158_n1681# a_n292_n1841# 1.75f
C5 a_n100_n1707# a_n292_n1841# 0.513f
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_F3SB2X a_n100_n1632# a_100_n1544# a_n292_n1766#
+ a_n158_n1544#
X0 a_100_n1544# a_n100_n1632# a_n158_n1544# a_n292_n1766# sky130_fd_pr__nfet_g5v0d10v5 ad=4.48 pd=31.5 as=4.48 ps=31.5 w=15.4 l=1
C0 a_n100_n1632# a_n158_n1544# 0.335f
C1 a_n100_n1632# a_100_n1544# 0.335f
C2 a_100_n1544# a_n158_n1544# 0.844f
C3 a_100_n1544# a_n292_n1766# 1.64f
C4 a_n158_n1544# a_n292_n1766# 1.64f
C5 a_n100_n1632# a_n292_n1766# 0.743f
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_2HXNYY a_n158_n1900# a_100_n1900# a_n292_n2122#
+ a_n100_n1988#
X0 a_100_n1900# a_n100_n1988# a_n158_n1900# a_n292_n2122# sky130_fd_pr__nfet_g5v0d10v5 ad=5.51 pd=38.6 as=5.51 ps=38.6 w=19 l=1
C0 a_n100_n1988# a_n158_n1900# 0.411f
C1 a_n100_n1988# a_100_n1900# 0.411f
C2 a_100_n1900# a_n158_n1900# 1.04f
C3 a_100_n1900# a_n292_n2122# 2.01f
C4 a_n158_n1900# a_n292_n2122# 2.01f
C5 a_n100_n1988# a_n292_n2122# 0.743f
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_24QKAW a_29_n1997# a_n487_n1997# a_487_n1900#
+ a_n287_n1900# a_n229_n1997# a_n545_n1900# a_n29_n1900# a_287_n1997# w_n745_n2197#
+ a_229_n1900# VSUBS
X0 a_487_n1900# a_287_n1997# a_229_n1900# w_n745_n2197# sky130_fd_pr__pfet_g5v0d10v5 ad=5.51 pd=38.6 as=2.76 ps=19.3 w=19 l=1
X1 a_n287_n1900# a_n487_n1997# a_n545_n1900# w_n745_n2197# sky130_fd_pr__pfet_g5v0d10v5 ad=2.76 pd=19.3 as=5.51 ps=38.6 w=19 l=1
X2 a_n29_n1900# a_n229_n1997# a_n287_n1900# w_n745_n2197# sky130_fd_pr__pfet_g5v0d10v5 ad=2.76 pd=19.3 as=2.76 ps=19.3 w=19 l=1
X3 a_229_n1900# a_29_n1997# a_n29_n1900# w_n745_n2197# sky130_fd_pr__pfet_g5v0d10v5 ad=2.76 pd=19.3 as=2.76 ps=19.3 w=19 l=1
C0 a_n287_n1900# a_n229_n1997# 0.411f
C1 w_n745_n2197# a_487_n1900# 1.09f
C2 w_n745_n2197# a_229_n1900# 0.022f
C3 w_n745_n2197# a_287_n1997# 0.386f
C4 a_n29_n1900# a_229_n1900# 1.04f
C5 w_n745_n2197# a_29_n1997# 0.343f
C6 a_n545_n1900# a_n287_n1900# 1.04f
C7 a_29_n1997# a_n29_n1900# 0.411f
C8 a_29_n1997# a_n229_n1997# 0.109f
C9 w_n745_n2197# a_n29_n1900# 0.022f
C10 w_n745_n2197# a_n487_n1997# 0.386f
C11 w_n745_n2197# a_n229_n1997# 0.343f
C12 a_n29_n1900# a_n229_n1997# 0.411f
C13 a_487_n1900# a_229_n1900# 1.04f
C14 a_n229_n1997# a_n487_n1997# 0.109f
C15 w_n745_n2197# a_n287_n1900# 0.022f
C16 w_n745_n2197# a_n545_n1900# 1.09f
C17 a_287_n1997# a_487_n1900# 0.411f
C18 a_n287_n1900# a_n29_n1900# 1.04f
C19 a_287_n1997# a_229_n1900# 0.411f
C20 a_29_n1997# a_229_n1900# 0.411f
C21 a_29_n1997# a_287_n1997# 0.109f
C22 a_n287_n1900# a_n487_n1997# 0.411f
C23 a_n545_n1900# a_n487_n1997# 0.411f
C24 a_487_n1900# VSUBS 0.925f
C25 a_229_n1900# VSUBS 0.527f
C26 a_n29_n1900# VSUBS 0.527f
C27 a_n287_n1900# VSUBS 0.527f
C28 a_n545_n1900# VSUBS 0.925f
C29 a_287_n1997# VSUBS 0.311f
C30 a_29_n1997# VSUBS 0.288f
C31 a_n229_n1997# VSUBS 0.288f
C32 a_n487_n1997# VSUBS 0.311f
C33 w_n745_n2197# VSUBS 22.5f
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_LB7Y8R a_n100_n157# a_n158_n69# a_n292_n291#
+ a_100_n69#
X0 a_100_n69# a_n100_n157# a_n158_n69# a_n292_n291# sky130_fd_pr__nfet_g5v0d10v5 ad=0.2 pd=1.96 as=0.2 ps=1.96 w=0.69 l=1
C0 a_n158_n69# a_100_n69# 0.0387f
C1 a_n100_n157# a_100_n69# 0.0202f
C2 a_n100_n157# a_n158_n69# 0.0202f
C3 a_100_n69# a_n292_n291# 0.105f
C4 a_n158_n69# a_n292_n291# 0.105f
C5 a_n100_n157# a_n292_n291# 0.683f
.ends

.subckt sky130_fd_pr__cap_mim_m3_1_8DB3RK m3_n876_n730# c1_n836_n690# VSUBS
X0 c1_n836_n690# m3_n876_n730# sky130_fd_pr__cap_mim_m3_1 l=6.9 w=6.9
C0 m3_n876_n730# c1_n836_n690# 4.73f
C1 c1_n836_n690# VSUBS 0.686f
C2 m3_n876_n730# VSUBS 2.42f
.ends

.subckt opamp VDD VSS V1 V2 VOUT
XXR3 VSS m1_4128_540# VOUT sky130_fd_pr__res_high_po_0p69_T8KQH6
XXM1 m1_5053_7611# VDD a_4864_8007# VDD VDD a_4864_8007# VSS sky130_fd_pr__pfet_g5v0d10v5_K8DQNF
XXM2 m1_4306_994# VSS V2 a_4864_8007# sky130_fd_pr__nfet_g5v0d10v5_VYCZE8
XXM3 a_4864_8007# VDD a_4864_8007# VDD VDD a_4864_8007# VSS sky130_fd_pr__pfet_g5v0d10v5_K8DQNF
XXM4 m1_5053_7611# VSS V1 m1_4306_994# sky130_fd_pr__nfet_g5v0d10v5_VYCZE8
XXM5 m1_5284_1188# VSS VSS m1_4306_994# sky130_fd_pr__nfet_g5v0d10v5_F3SB2X
XXM6 VSS VOUT VSS m1_5284_1188# sky130_fd_pr__nfet_g5v0d10v5_2HXNYY
XXM7 m1_5284_1188# m1_5284_1188# VSS VSS sky130_fd_pr__nfet_g5v0d10v5_F3SB2X
XXM8 m1_5053_7611# m1_5053_7611# VDD VOUT m1_5053_7611# VDD VDD m1_5053_7611# VDD
+ VOUT VSS sky130_fd_pr__pfet_g5v0d10v5_24QKAW
XXM9 VDD VDD VSS m1_5284_1188# sky130_fd_pr__nfet_g5v0d10v5_LB7Y8R
XXC1 m1_5053_7611# m1_4128_540# VSS sky130_fd_pr__cap_mim_m3_1_8DB3RK
C0 V1 m3_5211_1261# 0.14f
C1 m3_5211_1261# a_4864_8007# 0.0192f
C2 m3_5211_1261# VOUT 0.00865f
C3 m1_5284_1188# m1_4306_994# 2.09f
C4 m1_4306_994# VDD 0.00701f
C5 m1_4306_994# m1_4128_540# 0.354f
C6 m1_5284_1188# VDD 1.67f
C7 m1_5284_1188# m1_4128_540# 0.031f
C8 VDD m1_4128_540# 0.376f
C9 m1_4306_994# m1_5053_7611# 0.673f
C10 m1_5284_1188# m1_5053_7611# 0.0361f
C11 m1_5053_7611# VDD 10.4f
C12 m1_5053_7611# m1_4128_540# 0.115f
C13 m1_4306_994# V1 0.399f
C14 m3_5211_1261# V2 0.0767f
C15 m1_4306_994# a_4864_8007# 0.127f
C16 m1_5284_1188# V1 0.00363f
C17 V1 VDD 0.275f
C18 m1_4306_994# VOUT 0.00433f
C19 V1 m1_4128_540# 0.088f
C20 m1_5284_1188# a_4864_8007# 0.00623f
C21 VDD a_4864_8007# 1.96f
C22 m1_5284_1188# VOUT 2.28f
C23 VDD VOUT -1.29f
C24 a_4864_8007# m1_4128_540# 0.503f
C25 m1_4128_540# VOUT 0.00888f
C26 m1_5053_7611# V1 0.143f
C27 m1_5053_7611# a_4864_8007# 1.78f
C28 m1_5053_7611# VOUT 7.29f
C29 V1 a_4864_8007# 0.283f
C30 V1 VOUT 2.75e-19
C31 m1_4306_994# V2 0.213f
C32 a_4864_8007# VOUT 0.00842f
C33 m1_5284_1188# V2 9.56e-20
C34 VDD V2 0.00314f
C35 V2 m1_4128_540# 0.179f
C36 m1_4306_994# m3_5211_1261# 0.771f
C37 VDD m3_5211_1261# 0.0192f
C38 m1_5284_1188# m3_5211_1261# 0.446f
C39 m3_5211_1261# m1_4128_540# 0.0111f
C40 m1_5053_7611# V2 4.01e-19
C41 m1_5053_7611# m3_5211_1261# 0.0415f
C42 V1 V2 0.16f
C43 a_4864_8007# V2 0.263f
C44 m3_5211_1261# VSS 1.23f **FLOATING
C45 VDD VSS 46.6f
C46 m1_5053_7611# VSS 4.65f
C47 VOUT VSS 4.32f
C48 m1_5284_1188# VSS 8.17f
C49 V1 VSS 0.865f
C50 m1_4306_994# VSS 5.55f
C51 V2 VSS 0.848f
C52 a_4864_8007# VSS 4.88f
C53 m1_4128_540# VSS 2.47f
.ends

