magic
tech sky130A
magscale 1 2
timestamp 1720214482
<< nwell >>
rect -1777 -1797 1777 1797
<< mvpmos >>
rect -1519 -1500 -1319 1500
rect -1261 -1500 -1061 1500
rect -1003 -1500 -803 1500
rect -745 -1500 -545 1500
rect -487 -1500 -287 1500
rect -229 -1500 -29 1500
rect 29 -1500 229 1500
rect 287 -1500 487 1500
rect 545 -1500 745 1500
rect 803 -1500 1003 1500
rect 1061 -1500 1261 1500
rect 1319 -1500 1519 1500
<< mvpdiff >>
rect -1577 1488 -1519 1500
rect -1577 -1488 -1565 1488
rect -1531 -1488 -1519 1488
rect -1577 -1500 -1519 -1488
rect -1319 1488 -1261 1500
rect -1319 -1488 -1307 1488
rect -1273 -1488 -1261 1488
rect -1319 -1500 -1261 -1488
rect -1061 1488 -1003 1500
rect -1061 -1488 -1049 1488
rect -1015 -1488 -1003 1488
rect -1061 -1500 -1003 -1488
rect -803 1488 -745 1500
rect -803 -1488 -791 1488
rect -757 -1488 -745 1488
rect -803 -1500 -745 -1488
rect -545 1488 -487 1500
rect -545 -1488 -533 1488
rect -499 -1488 -487 1488
rect -545 -1500 -487 -1488
rect -287 1488 -229 1500
rect -287 -1488 -275 1488
rect -241 -1488 -229 1488
rect -287 -1500 -229 -1488
rect -29 1488 29 1500
rect -29 -1488 -17 1488
rect 17 -1488 29 1488
rect -29 -1500 29 -1488
rect 229 1488 287 1500
rect 229 -1488 241 1488
rect 275 -1488 287 1488
rect 229 -1500 287 -1488
rect 487 1488 545 1500
rect 487 -1488 499 1488
rect 533 -1488 545 1488
rect 487 -1500 545 -1488
rect 745 1488 803 1500
rect 745 -1488 757 1488
rect 791 -1488 803 1488
rect 745 -1500 803 -1488
rect 1003 1488 1061 1500
rect 1003 -1488 1015 1488
rect 1049 -1488 1061 1488
rect 1003 -1500 1061 -1488
rect 1261 1488 1319 1500
rect 1261 -1488 1273 1488
rect 1307 -1488 1319 1488
rect 1261 -1500 1319 -1488
rect 1519 1488 1577 1500
rect 1519 -1488 1531 1488
rect 1565 -1488 1577 1488
rect 1519 -1500 1577 -1488
<< mvpdiffc >>
rect -1565 -1488 -1531 1488
rect -1307 -1488 -1273 1488
rect -1049 -1488 -1015 1488
rect -791 -1488 -757 1488
rect -533 -1488 -499 1488
rect -275 -1488 -241 1488
rect -17 -1488 17 1488
rect 241 -1488 275 1488
rect 499 -1488 533 1488
rect 757 -1488 791 1488
rect 1015 -1488 1049 1488
rect 1273 -1488 1307 1488
rect 1531 -1488 1565 1488
<< mvnsubdiff >>
rect -1711 1719 1711 1731
rect -1711 1685 -1603 1719
rect 1603 1685 1711 1719
rect -1711 1673 1711 1685
rect -1711 1623 -1653 1673
rect -1711 -1623 -1699 1623
rect -1665 -1623 -1653 1623
rect 1653 1623 1711 1673
rect -1711 -1673 -1653 -1623
rect 1653 -1623 1665 1623
rect 1699 -1623 1711 1623
rect 1653 -1673 1711 -1623
rect -1711 -1685 1711 -1673
rect -1711 -1719 -1603 -1685
rect 1603 -1719 1711 -1685
rect -1711 -1731 1711 -1719
<< mvnsubdiffcont >>
rect -1603 1685 1603 1719
rect -1699 -1623 -1665 1623
rect 1665 -1623 1699 1623
rect -1603 -1719 1603 -1685
<< poly >>
rect -1519 1581 -1319 1597
rect -1519 1547 -1503 1581
rect -1335 1547 -1319 1581
rect -1519 1500 -1319 1547
rect -1261 1581 -1061 1597
rect -1261 1547 -1245 1581
rect -1077 1547 -1061 1581
rect -1261 1500 -1061 1547
rect -1003 1581 -803 1597
rect -1003 1547 -987 1581
rect -819 1547 -803 1581
rect -1003 1500 -803 1547
rect -745 1581 -545 1597
rect -745 1547 -729 1581
rect -561 1547 -545 1581
rect -745 1500 -545 1547
rect -487 1581 -287 1597
rect -487 1547 -471 1581
rect -303 1547 -287 1581
rect -487 1500 -287 1547
rect -229 1581 -29 1597
rect -229 1547 -213 1581
rect -45 1547 -29 1581
rect -229 1500 -29 1547
rect 29 1581 229 1597
rect 29 1547 45 1581
rect 213 1547 229 1581
rect 29 1500 229 1547
rect 287 1581 487 1597
rect 287 1547 303 1581
rect 471 1547 487 1581
rect 287 1500 487 1547
rect 545 1581 745 1597
rect 545 1547 561 1581
rect 729 1547 745 1581
rect 545 1500 745 1547
rect 803 1581 1003 1597
rect 803 1547 819 1581
rect 987 1547 1003 1581
rect 803 1500 1003 1547
rect 1061 1581 1261 1597
rect 1061 1547 1077 1581
rect 1245 1547 1261 1581
rect 1061 1500 1261 1547
rect 1319 1581 1519 1597
rect 1319 1547 1335 1581
rect 1503 1547 1519 1581
rect 1319 1500 1519 1547
rect -1519 -1547 -1319 -1500
rect -1519 -1581 -1503 -1547
rect -1335 -1581 -1319 -1547
rect -1519 -1597 -1319 -1581
rect -1261 -1547 -1061 -1500
rect -1261 -1581 -1245 -1547
rect -1077 -1581 -1061 -1547
rect -1261 -1597 -1061 -1581
rect -1003 -1547 -803 -1500
rect -1003 -1581 -987 -1547
rect -819 -1581 -803 -1547
rect -1003 -1597 -803 -1581
rect -745 -1547 -545 -1500
rect -745 -1581 -729 -1547
rect -561 -1581 -545 -1547
rect -745 -1597 -545 -1581
rect -487 -1547 -287 -1500
rect -487 -1581 -471 -1547
rect -303 -1581 -287 -1547
rect -487 -1597 -287 -1581
rect -229 -1547 -29 -1500
rect -229 -1581 -213 -1547
rect -45 -1581 -29 -1547
rect -229 -1597 -29 -1581
rect 29 -1547 229 -1500
rect 29 -1581 45 -1547
rect 213 -1581 229 -1547
rect 29 -1597 229 -1581
rect 287 -1547 487 -1500
rect 287 -1581 303 -1547
rect 471 -1581 487 -1547
rect 287 -1597 487 -1581
rect 545 -1547 745 -1500
rect 545 -1581 561 -1547
rect 729 -1581 745 -1547
rect 545 -1597 745 -1581
rect 803 -1547 1003 -1500
rect 803 -1581 819 -1547
rect 987 -1581 1003 -1547
rect 803 -1597 1003 -1581
rect 1061 -1547 1261 -1500
rect 1061 -1581 1077 -1547
rect 1245 -1581 1261 -1547
rect 1061 -1597 1261 -1581
rect 1319 -1547 1519 -1500
rect 1319 -1581 1335 -1547
rect 1503 -1581 1519 -1547
rect 1319 -1597 1519 -1581
<< polycont >>
rect -1503 1547 -1335 1581
rect -1245 1547 -1077 1581
rect -987 1547 -819 1581
rect -729 1547 -561 1581
rect -471 1547 -303 1581
rect -213 1547 -45 1581
rect 45 1547 213 1581
rect 303 1547 471 1581
rect 561 1547 729 1581
rect 819 1547 987 1581
rect 1077 1547 1245 1581
rect 1335 1547 1503 1581
rect -1503 -1581 -1335 -1547
rect -1245 -1581 -1077 -1547
rect -987 -1581 -819 -1547
rect -729 -1581 -561 -1547
rect -471 -1581 -303 -1547
rect -213 -1581 -45 -1547
rect 45 -1581 213 -1547
rect 303 -1581 471 -1547
rect 561 -1581 729 -1547
rect 819 -1581 987 -1547
rect 1077 -1581 1245 -1547
rect 1335 -1581 1503 -1547
<< locali >>
rect -1699 1685 -1603 1719
rect 1603 1685 1699 1719
rect -1699 1623 -1665 1685
rect 1665 1623 1699 1685
rect -1519 1547 -1503 1581
rect -1335 1547 -1319 1581
rect -1261 1547 -1245 1581
rect -1077 1547 -1061 1581
rect -1003 1547 -987 1581
rect -819 1547 -803 1581
rect -745 1547 -729 1581
rect -561 1547 -545 1581
rect -487 1547 -471 1581
rect -303 1547 -287 1581
rect -229 1547 -213 1581
rect -45 1547 -29 1581
rect 29 1547 45 1581
rect 213 1547 229 1581
rect 287 1547 303 1581
rect 471 1547 487 1581
rect 545 1547 561 1581
rect 729 1547 745 1581
rect 803 1547 819 1581
rect 987 1547 1003 1581
rect 1061 1547 1077 1581
rect 1245 1547 1261 1581
rect 1319 1547 1335 1581
rect 1503 1547 1519 1581
rect -1565 1488 -1531 1504
rect -1565 -1504 -1531 -1488
rect -1307 1488 -1273 1504
rect -1307 -1504 -1273 -1488
rect -1049 1488 -1015 1504
rect -1049 -1504 -1015 -1488
rect -791 1488 -757 1504
rect -791 -1504 -757 -1488
rect -533 1488 -499 1504
rect -533 -1504 -499 -1488
rect -275 1488 -241 1504
rect -275 -1504 -241 -1488
rect -17 1488 17 1504
rect -17 -1504 17 -1488
rect 241 1488 275 1504
rect 241 -1504 275 -1488
rect 499 1488 533 1504
rect 499 -1504 533 -1488
rect 757 1488 791 1504
rect 757 -1504 791 -1488
rect 1015 1488 1049 1504
rect 1015 -1504 1049 -1488
rect 1273 1488 1307 1504
rect 1273 -1504 1307 -1488
rect 1531 1488 1565 1504
rect 1531 -1504 1565 -1488
rect -1519 -1581 -1503 -1547
rect -1335 -1581 -1319 -1547
rect -1261 -1581 -1245 -1547
rect -1077 -1581 -1061 -1547
rect -1003 -1581 -987 -1547
rect -819 -1581 -803 -1547
rect -745 -1581 -729 -1547
rect -561 -1581 -545 -1547
rect -487 -1581 -471 -1547
rect -303 -1581 -287 -1547
rect -229 -1581 -213 -1547
rect -45 -1581 -29 -1547
rect 29 -1581 45 -1547
rect 213 -1581 229 -1547
rect 287 -1581 303 -1547
rect 471 -1581 487 -1547
rect 545 -1581 561 -1547
rect 729 -1581 745 -1547
rect 803 -1581 819 -1547
rect 987 -1581 1003 -1547
rect 1061 -1581 1077 -1547
rect 1245 -1581 1261 -1547
rect 1319 -1581 1335 -1547
rect 1503 -1581 1519 -1547
rect -1699 -1685 -1665 -1623
rect 1665 -1685 1699 -1623
rect -1699 -1719 -1603 -1685
rect 1603 -1719 1699 -1685
<< viali >>
rect -1503 1547 -1335 1581
rect -1245 1547 -1077 1581
rect -987 1547 -819 1581
rect -729 1547 -561 1581
rect -471 1547 -303 1581
rect -213 1547 -45 1581
rect 45 1547 213 1581
rect 303 1547 471 1581
rect 561 1547 729 1581
rect 819 1547 987 1581
rect 1077 1547 1245 1581
rect 1335 1547 1503 1581
rect -1565 -1488 -1531 1488
rect -1307 -1488 -1273 1488
rect -1049 -1488 -1015 1488
rect -791 -1488 -757 1488
rect -533 -1488 -499 1488
rect -275 -1488 -241 1488
rect -17 -1488 17 1488
rect 241 -1488 275 1488
rect 499 -1488 533 1488
rect 757 -1488 791 1488
rect 1015 -1488 1049 1488
rect 1273 -1488 1307 1488
rect 1531 -1488 1565 1488
rect -1503 -1581 -1335 -1547
rect -1245 -1581 -1077 -1547
rect -987 -1581 -819 -1547
rect -729 -1581 -561 -1547
rect -471 -1581 -303 -1547
rect -213 -1581 -45 -1547
rect 45 -1581 213 -1547
rect 303 -1581 471 -1547
rect 561 -1581 729 -1547
rect 819 -1581 987 -1547
rect 1077 -1581 1245 -1547
rect 1335 -1581 1503 -1547
<< metal1 >>
rect -1515 1581 -1323 1587
rect -1515 1547 -1503 1581
rect -1335 1547 -1323 1581
rect -1515 1541 -1323 1547
rect -1257 1581 -1065 1587
rect -1257 1547 -1245 1581
rect -1077 1547 -1065 1581
rect -1257 1541 -1065 1547
rect -999 1581 -807 1587
rect -999 1547 -987 1581
rect -819 1547 -807 1581
rect -999 1541 -807 1547
rect -741 1581 -549 1587
rect -741 1547 -729 1581
rect -561 1547 -549 1581
rect -741 1541 -549 1547
rect -483 1581 -291 1587
rect -483 1547 -471 1581
rect -303 1547 -291 1581
rect -483 1541 -291 1547
rect -225 1581 -33 1587
rect -225 1547 -213 1581
rect -45 1547 -33 1581
rect -225 1541 -33 1547
rect 33 1581 225 1587
rect 33 1547 45 1581
rect 213 1547 225 1581
rect 33 1541 225 1547
rect 291 1581 483 1587
rect 291 1547 303 1581
rect 471 1547 483 1581
rect 291 1541 483 1547
rect 549 1581 741 1587
rect 549 1547 561 1581
rect 729 1547 741 1581
rect 549 1541 741 1547
rect 807 1581 999 1587
rect 807 1547 819 1581
rect 987 1547 999 1581
rect 807 1541 999 1547
rect 1065 1581 1257 1587
rect 1065 1547 1077 1581
rect 1245 1547 1257 1581
rect 1065 1541 1257 1547
rect 1323 1581 1515 1587
rect 1323 1547 1335 1581
rect 1503 1547 1515 1581
rect 1323 1541 1515 1547
rect -1571 1488 -1525 1500
rect -1571 -1488 -1565 1488
rect -1531 -1488 -1525 1488
rect -1571 -1500 -1525 -1488
rect -1313 1488 -1267 1500
rect -1313 -1488 -1307 1488
rect -1273 -1488 -1267 1488
rect -1313 -1500 -1267 -1488
rect -1055 1488 -1009 1500
rect -1055 -1488 -1049 1488
rect -1015 -1488 -1009 1488
rect -1055 -1500 -1009 -1488
rect -797 1488 -751 1500
rect -797 -1488 -791 1488
rect -757 -1488 -751 1488
rect -797 -1500 -751 -1488
rect -539 1488 -493 1500
rect -539 -1488 -533 1488
rect -499 -1488 -493 1488
rect -539 -1500 -493 -1488
rect -281 1488 -235 1500
rect -281 -1488 -275 1488
rect -241 -1488 -235 1488
rect -281 -1500 -235 -1488
rect -23 1488 23 1500
rect -23 -1488 -17 1488
rect 17 -1488 23 1488
rect -23 -1500 23 -1488
rect 235 1488 281 1500
rect 235 -1488 241 1488
rect 275 -1488 281 1488
rect 235 -1500 281 -1488
rect 493 1488 539 1500
rect 493 -1488 499 1488
rect 533 -1488 539 1488
rect 493 -1500 539 -1488
rect 751 1488 797 1500
rect 751 -1488 757 1488
rect 791 -1488 797 1488
rect 751 -1500 797 -1488
rect 1009 1488 1055 1500
rect 1009 -1488 1015 1488
rect 1049 -1488 1055 1488
rect 1009 -1500 1055 -1488
rect 1267 1488 1313 1500
rect 1267 -1488 1273 1488
rect 1307 -1488 1313 1488
rect 1267 -1500 1313 -1488
rect 1525 1488 1571 1500
rect 1525 -1488 1531 1488
rect 1565 -1488 1571 1488
rect 1525 -1500 1571 -1488
rect -1515 -1547 -1323 -1541
rect -1515 -1581 -1503 -1547
rect -1335 -1581 -1323 -1547
rect -1515 -1587 -1323 -1581
rect -1257 -1547 -1065 -1541
rect -1257 -1581 -1245 -1547
rect -1077 -1581 -1065 -1547
rect -1257 -1587 -1065 -1581
rect -999 -1547 -807 -1541
rect -999 -1581 -987 -1547
rect -819 -1581 -807 -1547
rect -999 -1587 -807 -1581
rect -741 -1547 -549 -1541
rect -741 -1581 -729 -1547
rect -561 -1581 -549 -1547
rect -741 -1587 -549 -1581
rect -483 -1547 -291 -1541
rect -483 -1581 -471 -1547
rect -303 -1581 -291 -1547
rect -483 -1587 -291 -1581
rect -225 -1547 -33 -1541
rect -225 -1581 -213 -1547
rect -45 -1581 -33 -1547
rect -225 -1587 -33 -1581
rect 33 -1547 225 -1541
rect 33 -1581 45 -1547
rect 213 -1581 225 -1547
rect 33 -1587 225 -1581
rect 291 -1547 483 -1541
rect 291 -1581 303 -1547
rect 471 -1581 483 -1547
rect 291 -1587 483 -1581
rect 549 -1547 741 -1541
rect 549 -1581 561 -1547
rect 729 -1581 741 -1547
rect 549 -1587 741 -1581
rect 807 -1547 999 -1541
rect 807 -1581 819 -1547
rect 987 -1581 999 -1547
rect 807 -1587 999 -1581
rect 1065 -1547 1257 -1541
rect 1065 -1581 1077 -1547
rect 1245 -1581 1257 -1547
rect 1065 -1587 1257 -1581
rect 1323 -1547 1515 -1541
rect 1323 -1581 1335 -1547
rect 1503 -1581 1515 -1547
rect 1323 -1587 1515 -1581
<< properties >>
string FIXED_BBOX -1682 -1702 1682 1702
string gencell sky130_fd_pr__pfet_g5v0d10v5
string library sky130
string parameters w 15 l 1 m 1 nf 12 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
