magic
tech sky130A
timestamp 1716807968
<< pwell >>
rect -164 -329 164 329
<< mvnmos >>
rect -50 -200 50 200
<< mvndiff >>
rect -79 194 -50 200
rect -79 -194 -73 194
rect -56 -194 -50 194
rect -79 -200 -50 -194
rect 50 194 79 200
rect 50 -194 56 194
rect 73 -194 79 194
rect 50 -200 79 -194
<< mvndiffc >>
rect -73 -194 -56 194
rect 56 -194 73 194
<< mvpsubdiff >>
rect -146 305 146 311
rect -146 288 -92 305
rect 92 288 146 305
rect -146 282 146 288
rect -146 257 -117 282
rect -146 -257 -140 257
rect -123 -257 -117 257
rect 117 257 146 282
rect -146 -282 -117 -257
rect 117 -257 123 257
rect 140 -257 146 257
rect 117 -282 146 -257
rect -146 -288 146 -282
rect -146 -305 -92 -288
rect 92 -305 146 -288
rect -146 -311 146 -305
<< mvpsubdiffcont >>
rect -92 288 92 305
rect -140 -257 -123 257
rect 123 -257 140 257
rect -92 -305 92 -288
<< poly >>
rect -50 236 50 244
rect -50 219 -42 236
rect 42 219 50 236
rect -50 200 50 219
rect -50 -219 50 -200
rect -50 -236 -42 -219
rect 42 -236 50 -219
rect -50 -244 50 -236
<< polycont >>
rect -42 219 42 236
rect -42 -236 42 -219
<< locali >>
rect -140 288 -92 305
rect 92 288 140 305
rect -140 257 -123 288
rect 123 257 140 288
rect -50 219 -42 236
rect 42 219 50 236
rect -73 194 -56 202
rect -73 -202 -56 -194
rect 56 194 73 202
rect 56 -202 73 -194
rect -50 -236 -42 -219
rect 42 -236 50 -219
rect -140 -288 -123 -257
rect 123 -288 140 -257
rect -140 -305 -92 -288
rect 92 -305 140 -288
<< viali >>
rect -42 219 42 236
rect -73 -194 -56 194
rect 56 -194 73 194
rect -42 -236 42 -219
<< metal1 >>
rect -48 236 48 239
rect -48 219 -42 236
rect 42 219 48 236
rect -48 216 48 219
rect -76 194 -53 200
rect -76 -194 -73 194
rect -56 -194 -53 194
rect -76 -200 -53 -194
rect 53 194 76 200
rect 53 -194 56 194
rect 73 -194 76 194
rect 53 -200 76 -194
rect -48 -219 48 -216
rect -48 -236 -42 -219
rect 42 -236 48 -219
rect -48 -239 48 -236
<< properties >>
string FIXED_BBOX -131 -296 131 296
string gencell sky130_fd_pr__nfet_g5v0d10v5
string library sky130
string parameters w 4.0 l 1.0 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
