magic
tech sky130A
magscale 1 2
timestamp 1718246682
<< pwell >>
rect -586 -1804 586 1804
<< psubdiff >>
rect -550 1734 -454 1768
rect 454 1734 550 1768
rect -550 1672 -516 1734
rect 516 1672 550 1734
rect -550 -1734 -516 -1672
rect 516 -1734 550 -1672
rect -550 -1768 -454 -1734
rect 454 -1768 550 -1734
<< psubdiffcont >>
rect -454 1734 454 1768
rect -550 -1672 -516 1672
rect 516 -1672 550 1672
rect -454 -1768 454 -1734
<< xpolycontact >>
rect -420 1206 -282 1638
rect -420 -1638 -282 -1206
rect -186 1206 -48 1638
rect -186 -1638 -48 -1206
rect 48 1206 186 1638
rect 48 -1638 186 -1206
rect 282 1206 420 1638
rect 282 -1638 420 -1206
<< ppolyres >>
rect -420 -1206 -282 1206
rect -186 -1206 -48 1206
rect 48 -1206 186 1206
rect 282 -1206 420 1206
<< locali >>
rect -550 1734 -454 1768
rect 454 1734 550 1768
rect -550 1672 -516 1734
rect 516 1672 550 1734
rect -550 -1734 -516 -1672
rect 516 -1734 550 -1672
rect -550 -1768 -454 -1734
rect 454 -1768 550 -1734
<< viali >>
rect -404 1223 -298 1620
rect -170 1223 -64 1620
rect 64 1223 170 1620
rect 298 1223 404 1620
rect -404 -1620 -298 -1223
rect -170 -1620 -64 -1223
rect 64 -1620 170 -1223
rect 298 -1620 404 -1223
<< metal1 >>
rect -410 1620 -292 1632
rect -410 1223 -404 1620
rect -298 1223 -292 1620
rect -410 1211 -292 1223
rect -176 1620 -58 1632
rect -176 1223 -170 1620
rect -64 1223 -58 1620
rect -176 1211 -58 1223
rect 58 1620 176 1632
rect 58 1223 64 1620
rect 170 1223 176 1620
rect 58 1211 176 1223
rect 292 1620 410 1632
rect 292 1223 298 1620
rect 404 1223 410 1620
rect 292 1211 410 1223
rect -410 -1223 -292 -1211
rect -410 -1620 -404 -1223
rect -298 -1620 -292 -1223
rect -410 -1632 -292 -1620
rect -176 -1223 -58 -1211
rect -176 -1620 -170 -1223
rect -64 -1620 -58 -1223
rect -176 -1632 -58 -1620
rect 58 -1223 176 -1211
rect 58 -1620 64 -1223
rect 170 -1620 176 -1223
rect 58 -1632 176 -1620
rect 292 -1223 410 -1211
rect 292 -1620 298 -1223
rect 404 -1620 410 -1223
rect 292 -1632 410 -1620
<< properties >>
string FIXED_BBOX -533 -1751 533 1751
string gencell sky130_fd_pr__res_high_po_0p69
string library sky130
string parameters w 0.690 l 12.22 m 1 nx 4 wmin 0.690 lmin 0.50 rho 319.8 val 6.228k dummy 0 dw 0.0 term 194.82 sterm 0.0 caplen 0 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_high_po_0p35  sky130_fd_pr__res_high_po_0p69 sky130_fd_pr__res_high_po_1p41  sky130_fd_pr__res_high_po_2p85 sky130_fd_pr__res_high_po_5p73} snake 0 full_metal 1 wmax 0.690 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
