magic
tech sky130A
magscale 1 2
timestamp 1716807968
<< pwell >>
rect -586 -6874 586 6874
<< psubdiff >>
rect -550 6804 -454 6838
rect 454 6804 550 6838
rect -550 6742 -516 6804
rect 516 6742 550 6804
rect -550 -6804 -516 -6742
rect 516 -6804 550 -6742
rect -550 -6838 -454 -6804
rect 454 -6838 550 -6804
<< psubdiffcont >>
rect -454 6804 454 6838
rect -550 -6742 -516 6742
rect 516 -6742 550 6742
rect -454 -6838 454 -6804
<< xpolycontact >>
rect -420 6276 -282 6708
rect -420 3432 -282 3864
rect -186 6276 -48 6708
rect -186 3432 -48 3864
rect 48 6276 186 6708
rect 48 3432 186 3864
rect 282 6276 420 6708
rect 282 3432 420 3864
rect -420 2896 -282 3328
rect -420 52 -282 484
rect -186 2896 -48 3328
rect -186 52 -48 484
rect 48 2896 186 3328
rect 48 52 186 484
rect 282 2896 420 3328
rect 282 52 420 484
rect -420 -484 -282 -52
rect -420 -3328 -282 -2896
rect -186 -484 -48 -52
rect -186 -3328 -48 -2896
rect 48 -484 186 -52
rect 48 -3328 186 -2896
rect 282 -484 420 -52
rect 282 -3328 420 -2896
rect -420 -3864 -282 -3432
rect -420 -6708 -282 -6276
rect -186 -3864 -48 -3432
rect -186 -6708 -48 -6276
rect 48 -3864 186 -3432
rect 48 -6708 186 -6276
rect 282 -3864 420 -3432
rect 282 -6708 420 -6276
<< ppolyres >>
rect -420 3864 -282 6276
rect -186 3864 -48 6276
rect 48 3864 186 6276
rect 282 3864 420 6276
rect -420 484 -282 2896
rect -186 484 -48 2896
rect 48 484 186 2896
rect 282 484 420 2896
rect -420 -2896 -282 -484
rect -186 -2896 -48 -484
rect 48 -2896 186 -484
rect 282 -2896 420 -484
rect -420 -6276 -282 -3864
rect -186 -6276 -48 -3864
rect 48 -6276 186 -3864
rect 282 -6276 420 -3864
<< locali >>
rect -550 6804 -454 6838
rect 454 6804 550 6838
rect -550 6742 -516 6804
rect 516 6742 550 6804
rect -550 -6804 -516 -6742
rect 516 -6804 550 -6742
rect -550 -6838 -454 -6804
rect 454 -6838 550 -6804
<< viali >>
rect -404 6293 -298 6690
rect -170 6293 -64 6690
rect 64 6293 170 6690
rect 298 6293 404 6690
rect -404 3450 -298 3847
rect -170 3450 -64 3847
rect 64 3450 170 3847
rect 298 3450 404 3847
rect -404 2913 -298 3310
rect -170 2913 -64 3310
rect 64 2913 170 3310
rect 298 2913 404 3310
rect -404 70 -298 467
rect -170 70 -64 467
rect 64 70 170 467
rect 298 70 404 467
rect -404 -467 -298 -70
rect -170 -467 -64 -70
rect 64 -467 170 -70
rect 298 -467 404 -70
rect -404 -3310 -298 -2913
rect -170 -3310 -64 -2913
rect 64 -3310 170 -2913
rect 298 -3310 404 -2913
rect -404 -3847 -298 -3450
rect -170 -3847 -64 -3450
rect 64 -3847 170 -3450
rect 298 -3847 404 -3450
rect -404 -6690 -298 -6293
rect -170 -6690 -64 -6293
rect 64 -6690 170 -6293
rect 298 -6690 404 -6293
<< metal1 >>
rect -410 6690 -292 6702
rect -410 6293 -404 6690
rect -298 6293 -292 6690
rect -410 6281 -292 6293
rect -176 6690 -58 6702
rect -176 6293 -170 6690
rect -64 6293 -58 6690
rect -176 6281 -58 6293
rect 58 6690 176 6702
rect 58 6293 64 6690
rect 170 6293 176 6690
rect 58 6281 176 6293
rect 292 6690 410 6702
rect 292 6293 298 6690
rect 404 6293 410 6690
rect 292 6281 410 6293
rect -410 3847 -292 3859
rect -410 3450 -404 3847
rect -298 3450 -292 3847
rect -410 3438 -292 3450
rect -176 3847 -58 3859
rect -176 3450 -170 3847
rect -64 3450 -58 3847
rect -176 3438 -58 3450
rect 58 3847 176 3859
rect 58 3450 64 3847
rect 170 3450 176 3847
rect 58 3438 176 3450
rect 292 3847 410 3859
rect 292 3450 298 3847
rect 404 3450 410 3847
rect 292 3438 410 3450
rect -410 3310 -292 3322
rect -410 2913 -404 3310
rect -298 2913 -292 3310
rect -410 2901 -292 2913
rect -176 3310 -58 3322
rect -176 2913 -170 3310
rect -64 2913 -58 3310
rect -176 2901 -58 2913
rect 58 3310 176 3322
rect 58 2913 64 3310
rect 170 2913 176 3310
rect 58 2901 176 2913
rect 292 3310 410 3322
rect 292 2913 298 3310
rect 404 2913 410 3310
rect 292 2901 410 2913
rect -410 467 -292 479
rect -410 70 -404 467
rect -298 70 -292 467
rect -410 58 -292 70
rect -176 467 -58 479
rect -176 70 -170 467
rect -64 70 -58 467
rect -176 58 -58 70
rect 58 467 176 479
rect 58 70 64 467
rect 170 70 176 467
rect 58 58 176 70
rect 292 467 410 479
rect 292 70 298 467
rect 404 70 410 467
rect 292 58 410 70
rect -410 -70 -292 -58
rect -410 -467 -404 -70
rect -298 -467 -292 -70
rect -410 -479 -292 -467
rect -176 -70 -58 -58
rect -176 -467 -170 -70
rect -64 -467 -58 -70
rect -176 -479 -58 -467
rect 58 -70 176 -58
rect 58 -467 64 -70
rect 170 -467 176 -70
rect 58 -479 176 -467
rect 292 -70 410 -58
rect 292 -467 298 -70
rect 404 -467 410 -70
rect 292 -479 410 -467
rect -410 -2913 -292 -2901
rect -410 -3310 -404 -2913
rect -298 -3310 -292 -2913
rect -410 -3322 -292 -3310
rect -176 -2913 -58 -2901
rect -176 -3310 -170 -2913
rect -64 -3310 -58 -2913
rect -176 -3322 -58 -3310
rect 58 -2913 176 -2901
rect 58 -3310 64 -2913
rect 170 -3310 176 -2913
rect 58 -3322 176 -3310
rect 292 -2913 410 -2901
rect 292 -3310 298 -2913
rect 404 -3310 410 -2913
rect 292 -3322 410 -3310
rect -410 -3450 -292 -3438
rect -410 -3847 -404 -3450
rect -298 -3847 -292 -3450
rect -410 -3859 -292 -3847
rect -176 -3450 -58 -3438
rect -176 -3847 -170 -3450
rect -64 -3847 -58 -3450
rect -176 -3859 -58 -3847
rect 58 -3450 176 -3438
rect 58 -3847 64 -3450
rect 170 -3847 176 -3450
rect 58 -3859 176 -3847
rect 292 -3450 410 -3438
rect 292 -3847 298 -3450
rect 404 -3847 410 -3450
rect 292 -3859 410 -3847
rect -410 -6293 -292 -6281
rect -410 -6690 -404 -6293
rect -298 -6690 -292 -6293
rect -410 -6702 -292 -6690
rect -176 -6293 -58 -6281
rect -176 -6690 -170 -6293
rect -64 -6690 -58 -6293
rect -176 -6702 -58 -6690
rect 58 -6293 176 -6281
rect 58 -6690 64 -6293
rect 170 -6690 176 -6293
rect 58 -6702 176 -6690
rect 292 -6293 410 -6281
rect 292 -6690 298 -6293
rect 404 -6690 410 -6293
rect 292 -6702 410 -6690
<< properties >>
string FIXED_BBOX -533 -6821 533 6821
string gencell sky130_fd_pr__res_high_po_0p69
string library sky130
string parameters w 0.69 l 12.22 m 4 nx 4 wmin 0.690 lmin 0.50 rho 319.8 val 6.228k dummy 0 dw 0.0 term 194.82 sterm 0.0 caplen 0 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_high_po_0p35  sky130_fd_pr__res_high_po_0p69 sky130_fd_pr__res_high_po_1p41  sky130_fd_pr__res_high_po_2p85 sky130_fd_pr__res_high_po_5p73} snake 0 full_metal 1 wmax 0.690 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
