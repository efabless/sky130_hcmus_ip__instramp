magic
tech sky130A
magscale 1 2
timestamp 1716965124
<< pwell >>
rect 1828 -194 11784 4950
<< locali >>
rect 1906 1370 2004 4872
rect 2362 1370 2524 4872
rect 2890 1370 3168 4872
rect 1906 1364 3168 1370
rect 3758 1364 4090 4872
rect 1906 1354 4090 1364
rect 5160 1354 5538 4872
rect 7546 1354 7836 4872
rect 11712 1354 11736 4872
rect 1906 1248 11736 1354
rect 1906 1216 3088 1248
rect 3758 1246 11736 1248
rect 3882 1230 11736 1246
rect 2974 -124 3088 1216
rect 3872 1198 11736 1230
rect 3872 -124 3986 1198
rect 5284 1180 11736 1198
rect 5282 1154 11736 1180
rect 5282 -124 5396 1154
rect 7726 -124 7840 1154
<< metal1 >>
rect 2124 4395 11590 4736
rect 1690 4315 11590 4395
rect 2124 1470 2433 1893
rect 2651 1472 2960 1895
rect 1690 1072 2282 1202
rect 1690 1034 1990 1044
rect 1690 974 1920 1034
rect 1980 974 1990 1034
rect 1690 964 1990 974
rect 1690 926 1990 936
rect 1690 866 1920 926
rect 1980 866 1990 926
rect 1690 856 1990 866
rect 1690 818 1990 828
rect 1690 758 1920 818
rect 1980 758 1990 818
rect 1690 748 1990 758
rect 1690 710 1990 720
rect 1690 650 1920 710
rect 1980 650 1990 710
rect 1690 640 1990 650
rect 1690 603 1990 612
rect 1690 543 1920 603
rect 1980 543 1990 603
rect 1690 532 1990 543
rect 1690 376 2080 380
rect 1690 370 2089 376
rect 1690 310 2031 370
rect 2083 310 2089 370
rect 1690 304 2089 310
rect 1690 300 2080 304
rect 2120 31 2250 1072
rect 2315 896 2433 1470
rect 2646 1034 2776 1095
rect 2646 974 2681 1034
rect 2741 974 2776 1034
rect 2551 370 2615 376
rect 2551 310 2557 370
rect 2609 310 2615 370
rect 2551 304 2615 310
rect 2646 30 2776 974
rect 2842 896 2960 1472
rect 3284 1471 3844 1894
rect 4210 1472 5254 1894
rect 5664 1472 7704 1894
rect 3288 926 3418 1095
rect 3288 866 3330 926
rect 3390 866 3418 926
rect 3160 480 3240 490
rect 3160 420 3170 480
rect 3230 420 3240 480
rect 3160 410 3240 420
rect 3288 30 3418 866
rect 3544 926 3674 1095
rect 3544 866 3580 926
rect 3640 866 3674 926
rect 3447 370 3511 376
rect 3447 310 3453 370
rect 3505 310 3511 370
rect 3447 304 3511 310
rect 3544 30 3674 866
rect 3734 480 3843 1471
rect 4180 818 4310 1095
rect 4180 758 4220 818
rect 4280 758 4310 818
rect 3720 420 3730 480
rect 3830 420 3843 480
rect 3734 400 3843 420
rect 4060 480 4140 490
rect 4060 420 4068 480
rect 4130 420 4140 480
rect 4060 410 4140 420
rect 3734 344 3759 400
rect 4180 30 4310 758
rect 4440 818 4570 1095
rect 4440 758 4477 818
rect 4537 758 4570 818
rect 4343 370 4407 376
rect 4343 310 4349 370
rect 4401 310 4407 370
rect 4343 304 4407 310
rect 4440 30 4570 758
rect 4700 818 4830 1096
rect 4700 758 4736 818
rect 4796 758 4830 818
rect 4601 480 4665 486
rect 4601 420 4607 480
rect 4659 420 4665 480
rect 4601 414 4665 420
rect 4700 31 4830 758
rect 4958 818 5088 1096
rect 4958 758 4988 818
rect 5048 758 5088 818
rect 4859 370 4923 376
rect 4859 310 4865 370
rect 4917 310 4923 370
rect 4859 304 4923 310
rect 4958 31 5088 758
rect 5145 500 5254 1472
rect 5126 480 5254 500
rect 5596 710 5726 1095
rect 5596 650 5635 710
rect 5695 650 5726 710
rect 5126 420 5140 480
rect 5240 420 5254 480
rect 5126 400 5254 420
rect 5470 480 5552 490
rect 5470 420 5480 480
rect 5540 420 5552 480
rect 5470 410 5552 420
rect 5596 30 5726 650
rect 5855 710 5985 1096
rect 5855 650 5890 710
rect 5950 650 5985 710
rect 5755 370 5819 376
rect 5755 310 5761 370
rect 5813 310 5819 370
rect 5755 304 5819 310
rect 5855 31 5985 650
rect 6115 710 6245 1096
rect 6115 650 6150 710
rect 6210 650 6245 710
rect 6013 480 6077 490
rect 6013 420 6019 480
rect 6071 420 6077 480
rect 6013 410 6077 420
rect 6115 31 6245 650
rect 6373 710 6503 1096
rect 6373 650 6410 710
rect 6470 650 6503 710
rect 6273 370 6337 376
rect 6273 310 6278 370
rect 6330 310 6337 370
rect 6273 304 6337 310
rect 6373 31 6503 650
rect 6630 710 6760 1096
rect 6630 650 6665 710
rect 6725 650 6760 710
rect 6532 480 6596 490
rect 6532 420 6536 480
rect 6588 420 6596 480
rect 6532 410 6596 420
rect 6630 31 6760 650
rect 6887 710 7017 1096
rect 6887 650 6924 710
rect 6984 650 7017 710
rect 6789 370 6853 376
rect 6789 310 6793 370
rect 6845 310 6853 370
rect 6789 304 6853 310
rect 6887 31 7017 650
rect 7144 710 7274 1096
rect 7144 650 7180 710
rect 7240 650 7274 710
rect 7050 480 7114 490
rect 7050 420 7053 480
rect 7105 420 7114 480
rect 7050 410 7114 420
rect 7144 31 7274 650
rect 7400 710 7530 1096
rect 7400 650 7430 710
rect 7490 650 7530 710
rect 7304 370 7368 376
rect 7304 310 7310 370
rect 7362 310 7368 370
rect 7304 304 7368 310
rect 7400 31 7530 650
rect 7595 500 7704 1472
rect 7961 1471 11734 1894
rect 7570 480 7704 500
rect 8039 602 8169 1096
rect 8039 542 8078 602
rect 8138 542 8169 602
rect 7570 420 7590 480
rect 7690 420 7704 480
rect 7570 400 7704 420
rect 7940 480 8004 490
rect 7940 420 7946 480
rect 7998 420 8004 480
rect 7940 410 8004 420
rect 8039 31 8169 542
rect 8297 602 8427 1096
rect 8297 542 8340 602
rect 8400 542 8427 602
rect 8200 370 8264 376
rect 8200 310 8206 370
rect 8258 310 8264 370
rect 8200 304 8264 310
rect 8297 31 8427 542
rect 8556 602 8686 1096
rect 8556 542 8593 602
rect 8653 542 8686 602
rect 8457 480 8521 490
rect 8457 420 8463 480
rect 8515 420 8521 480
rect 8457 410 8521 420
rect 8556 31 8686 542
rect 8815 602 8945 1096
rect 8815 542 8855 602
rect 8915 542 8945 602
rect 8716 370 8780 376
rect 8716 310 8722 370
rect 8774 310 8780 370
rect 8716 304 8780 310
rect 8815 31 8945 542
rect 9070 602 9200 1096
rect 9070 542 9106 602
rect 9166 542 9200 602
rect 8973 480 9037 490
rect 8973 420 8979 480
rect 9031 420 9037 480
rect 8973 410 9037 420
rect 9070 31 9200 542
rect 9329 602 9459 1096
rect 9329 542 9366 602
rect 9426 542 9459 602
rect 9231 370 9295 376
rect 9231 310 9237 370
rect 9289 310 9295 370
rect 9231 304 9295 310
rect 9329 31 9459 542
rect 9588 602 9718 1096
rect 9588 542 9624 602
rect 9684 542 9718 602
rect 9489 480 9553 490
rect 9489 420 9495 480
rect 9547 420 9553 480
rect 9489 410 9553 420
rect 9588 31 9718 542
rect 9845 602 9975 1096
rect 9845 542 9880 602
rect 9940 542 9975 602
rect 9747 370 9811 376
rect 9747 310 9753 370
rect 9805 310 9811 370
rect 9747 304 9811 310
rect 9845 31 9975 542
rect 10104 602 10234 1096
rect 10104 542 10140 602
rect 10200 542 10234 602
rect 10005 480 10069 490
rect 10005 420 10011 480
rect 10063 420 10069 480
rect 10005 410 10069 420
rect 10104 31 10234 542
rect 10360 602 10490 1096
rect 10360 542 10395 602
rect 10455 542 10490 602
rect 10263 370 10327 376
rect 10263 310 10269 370
rect 10321 310 10327 370
rect 10263 304 10327 310
rect 10360 31 10490 542
rect 10620 602 10750 1096
rect 10620 542 10655 602
rect 10715 542 10750 602
rect 10521 480 10585 490
rect 10521 420 10527 480
rect 10579 420 10585 480
rect 10521 410 10585 420
rect 10620 31 10750 542
rect 10877 602 11007 1096
rect 10877 542 10915 602
rect 10975 542 11007 602
rect 10779 370 10843 376
rect 10779 310 10785 370
rect 10837 310 10843 370
rect 10779 304 10843 310
rect 10877 31 11007 542
rect 11135 602 11265 1096
rect 11135 542 11174 602
rect 11234 542 11265 602
rect 11038 480 11102 490
rect 11038 420 11044 480
rect 11096 420 11102 480
rect 11038 410 11102 420
rect 11135 31 11265 542
rect 11393 602 11523 1096
rect 11625 966 11734 1471
rect 11393 542 11420 602
rect 11480 542 11523 602
rect 11295 370 11359 376
rect 11295 310 11301 370
rect 11353 310 11359 370
rect 11295 304 11359 310
rect 11393 31 11523 542
rect 11586 490 11734 966
rect 11562 480 11734 490
rect 11562 420 11580 480
rect 11720 420 11734 480
rect 11562 410 11734 420
<< via1 >>
rect 1920 974 1980 1034
rect 1920 866 1980 926
rect 1920 758 1980 818
rect 1920 650 1980 710
rect 1920 543 1980 603
rect 2031 310 2083 370
rect 2681 974 2741 1034
rect 2557 310 2609 370
rect 3330 866 3390 926
rect 3170 420 3230 480
rect 3580 866 3640 926
rect 3453 310 3505 370
rect 4220 758 4280 818
rect 3730 420 3830 480
rect 4068 420 4128 480
rect 4477 758 4537 818
rect 4349 310 4401 370
rect 4736 758 4796 818
rect 4607 420 4659 480
rect 4988 758 5048 818
rect 4865 310 4917 370
rect 5635 650 5695 710
rect 5140 420 5240 480
rect 5480 420 5540 480
rect 5890 650 5950 710
rect 5761 310 5813 370
rect 6150 650 6210 710
rect 6019 420 6071 480
rect 6410 650 6470 710
rect 6278 310 6330 370
rect 6665 650 6725 710
rect 6536 420 6588 480
rect 6924 650 6984 710
rect 6793 310 6845 370
rect 7180 650 7240 710
rect 7053 420 7105 480
rect 7430 650 7490 710
rect 7310 310 7362 370
rect 8078 542 8138 602
rect 7590 420 7690 480
rect 7946 420 7998 480
rect 8340 542 8400 602
rect 8206 310 8258 370
rect 8593 542 8653 602
rect 8463 420 8515 480
rect 8855 542 8915 602
rect 8722 310 8774 370
rect 9106 542 9166 602
rect 8979 420 9031 480
rect 9366 542 9426 602
rect 9237 310 9289 370
rect 9624 542 9684 602
rect 9495 420 9547 480
rect 9880 542 9940 602
rect 9753 310 9805 370
rect 10140 542 10200 602
rect 10011 420 10063 480
rect 10395 542 10455 602
rect 10269 310 10321 370
rect 10655 542 10715 602
rect 10527 420 10579 480
rect 10915 542 10975 602
rect 10785 310 10837 370
rect 11174 542 11234 602
rect 11044 420 11096 480
rect 11420 542 11480 602
rect 11301 310 11353 370
rect 11580 420 11720 480
<< metal2 >>
rect 1920 1034 2741 1044
rect 1980 974 2681 1034
rect 1920 964 2741 974
rect 1920 926 3640 936
rect 1980 866 3330 926
rect 3390 866 3580 926
rect 1920 856 3640 866
rect 1920 818 5070 828
rect 1980 758 4220 818
rect 4280 758 4477 818
rect 4537 758 4736 818
rect 4796 758 4988 818
rect 5048 758 5070 818
rect 1920 748 5070 758
rect 1920 710 7510 720
rect 1980 650 5635 710
rect 5695 650 5890 710
rect 5950 650 6150 710
rect 6210 650 6410 710
rect 6470 650 6665 710
rect 6725 650 6924 710
rect 6984 650 7180 710
rect 7240 650 7430 710
rect 7490 650 7510 710
rect 1920 640 7510 650
rect 1920 603 11500 612
rect 1980 602 11500 603
rect 1980 543 8078 602
rect 1920 542 8078 543
rect 8138 542 8340 602
rect 8400 542 8593 602
rect 8653 542 8855 602
rect 8915 542 9106 602
rect 9166 542 9366 602
rect 9426 542 9624 602
rect 9684 542 9880 602
rect 9940 542 10140 602
rect 10200 542 10395 602
rect 10455 542 10655 602
rect 10715 542 10915 602
rect 10975 542 11174 602
rect 11234 542 11420 602
rect 11480 542 11500 602
rect 1920 532 11500 542
rect 3160 480 3830 490
rect 3160 420 3170 480
rect 3230 420 3730 480
rect 3160 410 3830 420
rect 4060 480 5240 490
rect 4060 420 4068 480
rect 4128 420 4607 480
rect 4659 420 5140 480
rect 4060 410 5240 420
rect 5470 480 7690 490
rect 5470 420 5480 480
rect 5540 420 6019 480
rect 6071 420 6536 480
rect 6588 420 7053 480
rect 7105 420 7590 480
rect 5470 410 7690 420
rect 7940 480 11734 490
rect 7940 420 7946 480
rect 7998 420 8463 480
rect 8515 420 8979 480
rect 9031 420 9495 480
rect 9547 420 10011 480
rect 10063 420 10527 480
rect 10579 420 11044 480
rect 11096 420 11580 480
rect 11720 420 11734 480
rect 7940 410 11734 420
rect 2025 370 11359 376
rect 2025 310 2031 370
rect 2083 310 2557 370
rect 2609 310 3453 370
rect 3505 310 4349 370
rect 4401 310 4865 370
rect 4917 310 5761 370
rect 5813 310 6278 370
rect 6330 310 6793 370
rect 6845 310 7310 370
rect 7362 310 8206 370
rect 8258 310 8722 370
rect 8774 310 9237 370
rect 9289 310 9753 370
rect 9805 310 10269 370
rect 10321 310 10785 370
rect 10837 310 11301 370
rect 11353 310 11359 370
rect 2025 304 11359 310
use sky130_fd_pr__nfet_g5v0d10v5_727CUP  XM6
timestamp 1716884908
transform 1 0 2712 0 1 563
box -328 -735 328 735
use sky130_fd_pr__nfet_g5v0d10v5_VU5C5A  XM7
timestamp 1716884908
transform 1 0 3479 0 1 573
box -457 -745 457 745
use sky130_fd_pr__nfet_g5v0d10v5_S7E57E  XM8
timestamp 1716884908
transform 1 0 4633 0 1 551
box -715 -723 715 723
use sky130_fd_pr__nfet_g5v0d10v5_J97EKB  XM9
timestamp 1716884908
transform 1 0 6561 0 1 524
box -1231 -696 1231 696
use sky130_fd_pr__nfet_g5v0d10v5_YPGNM4  XM10
timestamp 1716884908
transform 1 0 9779 0 1 526
box -2005 -698 2005 698
use sky130_fd_pr__nfet_g5v0d10v5_727CUP  XM11
timestamp 1716884908
transform 1 0 2186 0 1 563
box -328 -735 328 735
use sky130_fd_pr__res_high_po_0p69_JKKHRG  XR1
timestamp 1716884908
transform 1 0 2711 0 1 3104
box -235 -1804 235 1804
use sky130_fd_pr__res_high_po_0p69_JKKHRG  XR2
timestamp 1716884908
transform 1 0 2183 0 1 3104
box -235 -1804 235 1804
use sky130_fd_pr__res_high_po_0p69_Z3RMRJ  XR3
timestamp 1716884908
transform 1 0 3460 0 1 3104
box -352 -1804 352 1804
use sky130_fd_pr__res_high_po_0p69_YMHKRJ  XR4
timestamp 1716884908
transform 1 0 4620 0 1 3104
box -586 -1804 586 1804
use sky130_fd_pr__res_high_po_0p69_Z3RMR6  XR5
timestamp 1716884908
transform 1 0 6542 0 1 3104
box -1054 -1804 1054 1804
use sky130_fd_pr__res_high_po_0p69_HBQF5Z  XR6
timestamp 1716884908
transform 1 0 9776 0 1 3104
box -1990 -1804 1990 1804
<< labels >>
rlabel metal1 1690 1072 1810 1192 0 VDD
port 1 nsew
rlabel locali 1912 1222 2032 1342 0 VSS
port 2 nsew
rlabel metal1 1690 300 1770 380 0 R1
port 4 nsew
rlabel metal1 1690 964 1770 1044 0 D0
port 5 nsew
rlabel metal1 1690 856 1770 936 0 D1
port 6 nsew
rlabel metal1 1690 748 1770 828 0 D2
port 7 nsew
rlabel metal1 1690 640 1770 720 0 D3
port 8 nsew
rlabel metal1 1690 532 1770 612 0 D4
port 9 nsew
rlabel metal1 1690 4315 1770 4395 0 R2
port 3 nsew
<< end >>
