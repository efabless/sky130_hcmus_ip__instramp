magic
tech sky130A
magscale 1 2
timestamp 1716453420
<< nwell >>
rect -487 -1797 487 1797
<< mvpmos >>
rect -229 -1500 -29 1500
rect 29 -1500 229 1500
<< mvpdiff >>
rect -287 1488 -229 1500
rect -287 -1488 -275 1488
rect -241 -1488 -229 1488
rect -287 -1500 -229 -1488
rect -29 1488 29 1500
rect -29 -1488 -17 1488
rect 17 -1488 29 1488
rect -29 -1500 29 -1488
rect 229 1488 287 1500
rect 229 -1488 241 1488
rect 275 -1488 287 1488
rect 229 -1500 287 -1488
<< mvpdiffc >>
rect -275 -1488 -241 1488
rect -17 -1488 17 1488
rect 241 -1488 275 1488
<< mvnsubdiff >>
rect -421 1719 421 1731
rect -421 1685 -313 1719
rect 313 1685 421 1719
rect -421 1673 421 1685
rect -421 1623 -363 1673
rect -421 -1623 -409 1623
rect -375 -1623 -363 1623
rect 363 1623 421 1673
rect -421 -1673 -363 -1623
rect 363 -1623 375 1623
rect 409 -1623 421 1623
rect 363 -1673 421 -1623
rect -421 -1685 421 -1673
rect -421 -1719 -313 -1685
rect 313 -1719 421 -1685
rect -421 -1731 421 -1719
<< mvnsubdiffcont >>
rect -313 1685 313 1719
rect -409 -1623 -375 1623
rect 375 -1623 409 1623
rect -313 -1719 313 -1685
<< poly >>
rect -229 1581 -29 1597
rect -229 1547 -213 1581
rect -45 1547 -29 1581
rect -229 1500 -29 1547
rect 29 1581 229 1597
rect 29 1547 45 1581
rect 213 1547 229 1581
rect 29 1500 229 1547
rect -229 -1547 -29 -1500
rect -229 -1581 -213 -1547
rect -45 -1581 -29 -1547
rect -229 -1597 -29 -1581
rect 29 -1547 229 -1500
rect 29 -1581 45 -1547
rect 213 -1581 229 -1547
rect 29 -1597 229 -1581
<< polycont >>
rect -213 1547 -45 1581
rect 45 1547 213 1581
rect -213 -1581 -45 -1547
rect 45 -1581 213 -1547
<< locali >>
rect -409 1685 -313 1719
rect 313 1685 409 1719
rect -409 1623 -375 1685
rect 375 1623 409 1685
rect -229 1547 -213 1581
rect -45 1547 -29 1581
rect 29 1547 45 1581
rect 213 1547 229 1581
rect -275 1488 -241 1504
rect -275 -1504 -241 -1488
rect -17 1488 17 1504
rect -17 -1504 17 -1488
rect 241 1488 275 1504
rect 241 -1504 275 -1488
rect -229 -1581 -213 -1547
rect -45 -1581 -29 -1547
rect 29 -1581 45 -1547
rect 213 -1581 229 -1547
rect -409 -1685 -375 -1623
rect 375 -1685 409 -1623
rect -409 -1719 -313 -1685
rect 313 -1719 409 -1685
<< viali >>
rect -213 1547 -45 1581
rect 45 1547 213 1581
rect -275 -1488 -241 1488
rect -17 -1488 17 1488
rect 241 -1488 275 1488
rect -213 -1581 -45 -1547
rect 45 -1581 213 -1547
<< metal1 >>
rect -225 1581 -33 1587
rect -225 1547 -213 1581
rect -45 1547 -33 1581
rect -225 1541 -33 1547
rect 33 1581 225 1587
rect 33 1547 45 1581
rect 213 1547 225 1581
rect 33 1541 225 1547
rect -281 1488 -235 1500
rect -281 -1488 -275 1488
rect -241 -1488 -235 1488
rect -281 -1500 -235 -1488
rect -23 1488 23 1500
rect -23 -1488 -17 1488
rect 17 -1488 23 1488
rect -23 -1500 23 -1488
rect 235 1488 281 1500
rect 235 -1488 241 1488
rect 275 -1488 281 1488
rect 235 -1500 281 -1488
rect -225 -1547 -33 -1541
rect -225 -1581 -213 -1547
rect -45 -1581 -33 -1547
rect -225 -1587 -33 -1581
rect 33 -1547 225 -1541
rect 33 -1581 45 -1547
rect 213 -1581 225 -1547
rect 33 -1587 225 -1581
<< properties >>
string FIXED_BBOX -392 -1702 392 1702
string gencell sky130_fd_pr__pfet_g5v0d10v5
string library sky130
string parameters w 15.0 l 1.0 m 1 nf 2 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
